--------------------------------------------------------------------------------
-- $RCSfile: $
--
-- DESC    : OpenRisk 1420 
--
-- AUTHOR  : Dr. Theo Kluter
--
-- CVS     : $Revision: $
--           $Date: $
--           $Author: $
--           $Source: $
--
--------------------------------------------------------------------------------
--
--  HISTORY :
--
--  $Log: 
--------------------------------------------------------------------------------

ARCHITECTURE platform_independent OF bios_rom IS

BEGIN

   TheRom : PROCESS( address )
   BEGIN
      CASE (address) IS
         WHEN "000000000000" => data <= X"0013ADDE";
         WHEN "000000000001" => data <= X"00000015";
         WHEN "000000000010" => data <= X"21000000";
         WHEN "000000000011" => data <= X"00000015";
         WHEN "000000000100" => data <= X"1F000000";
         WHEN "000000000101" => data <= X"00000015";
         WHEN "000000000110" => data <= X"1D000000";
         WHEN "000000000111" => data <= X"00000015";
         WHEN "000000001000" => data <= X"1B000000";
         WHEN "000000001001" => data <= X"00000015";
         WHEN "000000001010" => data <= X"19000000";
         WHEN "000000001011" => data <= X"00000015";
         WHEN "000000001100" => data <= X"17000000";
         WHEN "000000001101" => data <= X"00000015";
         WHEN "000000001110" => data <= X"15000000";
         WHEN "000000001111" => data <= X"00000015";
         WHEN "000000010000" => data <= X"13000000";
         WHEN "000000010001" => data <= X"00000015";
         WHEN "000000010010" => data <= X"11000000";
         WHEN "000000010011" => data <= X"00000015";
         WHEN "000000010100" => data <= X"0F000000";
         WHEN "000000010101" => data <= X"00000015";
         WHEN "000000010110" => data <= X"0D000000";
         WHEN "000000010111" => data <= X"00000015";
         WHEN "000000011000" => data <= X"0B000000";
         WHEN "000000011001" => data <= X"00000015";
         WHEN "000000011010" => data <= X"09000000";
         WHEN "000000011011" => data <= X"00000015";
         WHEN "000000011100" => data <= X"00C02018";
         WHEN "000000011101" => data <= X"FC1F21A8";
         WHEN "000000011110" => data <= X"050060E0";
         WHEN "000000011111" => data <= X"4B030004";
         WHEN "000000100000" => data <= X"050080E0";
         WHEN "000000100010" => data <= X"00000015";
         WHEN "000000100011" => data <= X"84FF219C";
         WHEN "000000100100" => data <= X"001001D4";
         WHEN "000000100101" => data <= X"041801D4";
         WHEN "000000100110" => data <= X"082001D4";
         WHEN "000000100111" => data <= X"0C2801D4";
         WHEN "000000101000" => data <= X"103001D4";
         WHEN "000000101001" => data <= X"143801D4";
         WHEN "000000101010" => data <= X"184001D4";
         WHEN "000000101011" => data <= X"1C4801D4";
         WHEN "000000101100" => data <= X"205001D4";
         WHEN "000000101101" => data <= X"245801D4";
         WHEN "000000101110" => data <= X"286001D4";
         WHEN "000000101111" => data <= X"2C6801D4";
         WHEN "000000110000" => data <= X"307001D4";
         WHEN "000000110001" => data <= X"347801D4";
         WHEN "000000110010" => data <= X"388001D4";
         WHEN "000000110011" => data <= X"3C8801D4";
         WHEN "000000110100" => data <= X"409001D4";
         WHEN "000000110101" => data <= X"449801D4";
         WHEN "000000110110" => data <= X"48A001D4";
         WHEN "000000110111" => data <= X"4CA801D4";
         WHEN "000000111000" => data <= X"50B001D4";
         WHEN "000000111001" => data <= X"54B801D4";
         WHEN "000000111010" => data <= X"58C001D4";
         WHEN "000000111011" => data <= X"5CC801D4";
         WHEN "000000111100" => data <= X"60D001D4";
         WHEN "000000111101" => data <= X"64D801D4";
         WHEN "000000111110" => data <= X"68E001D4";
         WHEN "000000111111" => data <= X"6CE801D4";
         WHEN "000001000000" => data <= X"70F001D4";
         WHEN "000001000001" => data <= X"74F801D4";
         WHEN "000001000010" => data <= X"1200E0B7";
         WHEN "000001000011" => data <= X"0200FFBB";
         WHEN "000001000100" => data <= X"00F0C01B";
         WHEN "000001000101" => data <= X"AC01DEAB";
         WHEN "000001000110" => data <= X"00F8DEE3";
         WHEN "000001000111" => data <= X"0000FE87";
         WHEN "000001001000" => data <= X"00F80048";
         WHEN "000001001001" => data <= X"00000015";
         WHEN "000001001010" => data <= X"00004184";
         WHEN "000001001011" => data <= X"04006184";
         WHEN "000001001100" => data <= X"08008184";
         WHEN "000001001101" => data <= X"0C00A184";
         WHEN "000001001110" => data <= X"1000C184";
         WHEN "000001001111" => data <= X"1400E184";
         WHEN "000001010000" => data <= X"18000185";
         WHEN "000001010001" => data <= X"1C002185";
         WHEN "000001010010" => data <= X"20004185";
         WHEN "000001010011" => data <= X"24006185";
         WHEN "000001010100" => data <= X"28008185";
         WHEN "000001010101" => data <= X"2C00A185";
         WHEN "000001010110" => data <= X"3000C185";
         WHEN "000001010111" => data <= X"3400E185";
         WHEN "000001011000" => data <= X"38000186";
         WHEN "000001011001" => data <= X"3C002186";
         WHEN "000001011010" => data <= X"40004186";
         WHEN "000001011011" => data <= X"44006186";
         WHEN "000001011100" => data <= X"48008186";
         WHEN "000001011101" => data <= X"4C00A186";
         WHEN "000001011110" => data <= X"5000C186";
         WHEN "000001011111" => data <= X"5400E186";
         WHEN "000001100000" => data <= X"58000187";
         WHEN "000001100001" => data <= X"5C002187";
         WHEN "000001100010" => data <= X"60004187";
         WHEN "000001100011" => data <= X"64006187";
         WHEN "000001100100" => data <= X"68008187";
         WHEN "000001100101" => data <= X"6C00A187";
         WHEN "000001100110" => data <= X"7000C187";
         WHEN "000001100111" => data <= X"7400E187";
         WHEN "000001101000" => data <= X"7C00219C";
         WHEN "000001101001" => data <= X"00000024";
         WHEN "000001101010" => data <= X"00000015";
         WHEN "000001101011" => data <= X"700000F0";
         WHEN "000001101100" => data <= X"E40100F0";
         WHEN "000001101101" => data <= X"000200F0";
         WHEN "000001101110" => data <= X"1C0200F0";
         WHEN "000001101111" => data <= X"380200F0";
         WHEN "000001110000" => data <= X"540200F0";
         WHEN "000001110001" => data <= X"700200F0";
         WHEN "000001110010" => data <= X"8C0200F0";
         WHEN "000001110011" => data <= X"A80200F0";
         WHEN "000001110100" => data <= X"C40200F0";
         WHEN "000001110101" => data <= X"E00200F0";
         WHEN "000001110110" => data <= X"FC0200F0";
         WHEN "000001110111" => data <= X"340300F0";
         WHEN "000001111000" => data <= X"180300F0";
         WHEN "000001111001" => data <= X"00F0A018";
         WHEN "000001111010" => data <= X"00F08018";
         WHEN "000001111011" => data <= X"00F06018";
         WHEN "000001111100" => data <= X"C01AA59C";
         WHEN "000001111101" => data <= X"B009849C";
         WHEN "000001111110" => data <= X"6A010000";
         WHEN "000001111111" => data <= X"180B639C";
         WHEN "000010000000" => data <= X"00F0A018";
         WHEN "000010000001" => data <= X"00F08018";
         WHEN "000010000010" => data <= X"00F06018";
         WHEN "000010000011" => data <= X"CC1AA59C";
         WHEN "000010000100" => data <= X"B009849C";
         WHEN "000010000101" => data <= X"63010000";
         WHEN "000010000110" => data <= X"180B639C";
         WHEN "000010000111" => data <= X"00F0A018";
         WHEN "000010001000" => data <= X"00F08018";
         WHEN "000010001001" => data <= X"00F06018";
         WHEN "000010001010" => data <= X"DD1AA59C";
         WHEN "000010001011" => data <= X"B009849C";
         WHEN "000010001100" => data <= X"5C010000";
         WHEN "000010001101" => data <= X"180B639C";
         WHEN "000010001110" => data <= X"00F0A018";
         WHEN "000010001111" => data <= X"00F08018";
         WHEN "000010010000" => data <= X"00F06018";
         WHEN "000010010001" => data <= X"EB1AA59C";
         WHEN "000010010010" => data <= X"B009849C";
         WHEN "000010010011" => data <= X"55010000";
         WHEN "000010010100" => data <= X"180B639C";
         WHEN "000010010101" => data <= X"00F0A018";
         WHEN "000010010110" => data <= X"00F08018";
         WHEN "000010010111" => data <= X"00F06018";
         WHEN "000010011000" => data <= X"F11AA59C";
         WHEN "000010011001" => data <= X"B009849C";
         WHEN "000010011010" => data <= X"4E010000";
         WHEN "000010011011" => data <= X"180B639C";
         WHEN "000010011100" => data <= X"00F0A018";
         WHEN "000010011101" => data <= X"00F08018";
         WHEN "000010011110" => data <= X"00F06018";
         WHEN "000010011111" => data <= X"FA1AA59C";
         WHEN "000010100000" => data <= X"B009849C";
         WHEN "000010100001" => data <= X"47010000";
         WHEN "000010100010" => data <= X"180B639C";
         WHEN "000010100011" => data <= X"00F0A018";
         WHEN "000010100100" => data <= X"00F08018";
         WHEN "000010100101" => data <= X"00F06018";
         WHEN "000010100110" => data <= X"001BA59C";
         WHEN "000010100111" => data <= X"B009849C";
         WHEN "000010101000" => data <= X"40010000";
         WHEN "000010101001" => data <= X"180B639C";
         WHEN "000010101010" => data <= X"00F0A018";
         WHEN "000010101011" => data <= X"00F08018";
         WHEN "000010101100" => data <= X"00F06018";
         WHEN "000010101101" => data <= X"061BA59C";
         WHEN "000010101110" => data <= X"B009849C";
         WHEN "000010101111" => data <= X"39010000";
         WHEN "000010110000" => data <= X"180B639C";
         WHEN "000010110001" => data <= X"00F0A018";
         WHEN "000010110010" => data <= X"00F08018";
         WHEN "000010110011" => data <= X"00F06018";
         WHEN "000010110100" => data <= X"0C1BA59C";
         WHEN "000010110101" => data <= X"B009849C";
         WHEN "000010110110" => data <= X"32010000";
         WHEN "000010110111" => data <= X"180B639C";
         WHEN "000010111000" => data <= X"00F0A018";
         WHEN "000010111001" => data <= X"00F08018";
         WHEN "000010111010" => data <= X"00F06018";
         WHEN "000010111011" => data <= X"121BA59C";
         WHEN "000010111100" => data <= X"B009849C";
         WHEN "000010111101" => data <= X"2B010000";
         WHEN "000010111110" => data <= X"180B639C";
         WHEN "000010111111" => data <= X"00F0A018";
         WHEN "000011000000" => data <= X"00F08018";
         WHEN "000011000001" => data <= X"00F06018";
         WHEN "000011000010" => data <= X"1A1BA59C";
         WHEN "000011000011" => data <= X"B009849C";
         WHEN "000011000100" => data <= X"24010000";
         WHEN "000011000101" => data <= X"180B639C";
         WHEN "000011000110" => data <= X"00F0A018";
         WHEN "000011000111" => data <= X"00F08018";
         WHEN "000011001000" => data <= X"00F06018";
         WHEN "000011001001" => data <= X"231BA59C";
         WHEN "000011001010" => data <= X"B009849C";
         WHEN "000011001011" => data <= X"1D010000";
         WHEN "000011001100" => data <= X"180B639C";
         WHEN "000011001101" => data <= X"00F0A018";
         WHEN "000011001110" => data <= X"00F08018";
         WHEN "000011001111" => data <= X"00F06018";
         WHEN "000011010000" => data <= X"2A1BA59C";
         WHEN "000011010001" => data <= X"B009849C";
         WHEN "000011010010" => data <= X"16010000";
         WHEN "000011010011" => data <= X"180B639C";
         WHEN "000011010100" => data <= X"0000601A";
         WHEN "000011010101" => data <= X"0700A0AA";
         WHEN "000011010110" => data <= X"02A83372";
         WHEN "000011010111" => data <= X"0000E01A";
         WHEN "000011011000" => data <= X"010031A6";
         WHEN "000011011001" => data <= X"00B831E4";
         WHEN "000011011010" => data <= X"FCFFFF13";
         WHEN "000011011011" => data <= X"00000015";
         WHEN "000011011100" => data <= X"00480044";
         WHEN "000011011101" => data <= X"00000015";
         WHEN "000011011110" => data <= X"00006019";
         WHEN "000011011111" => data <= X"02186B71";
         WHEN "000011100000" => data <= X"00480044";
         WHEN "000011100001" => data <= X"00000015";
         WHEN "000011100010" => data <= X"160020AA";
         WHEN "000011100011" => data <= X"02890370";
         WHEN "000011100100" => data <= X"020020AA";
         WHEN "000011100101" => data <= X"070060AA";
         WHEN "000011100110" => data <= X"02991170";
         WHEN "000011100111" => data <= X"EDFFFF03";
         WHEN "000011101000" => data <= X"00000015";
         WHEN "000011101001" => data <= X"DCFF219C";
         WHEN "000011101010" => data <= X"008001D4";
         WHEN "000011101011" => data <= X"049001D4";
         WHEN "000011101100" => data <= X"08A001D4";
         WHEN "000011101101" => data <= X"0CB001D4";
         WHEN "000011101110" => data <= X"10C001D4";
         WHEN "000011101111" => data <= X"14D001D4";
         WHEN "000011110000" => data <= X"18E001D4";
         WHEN "000011110001" => data <= X"1CF001D4";
         WHEN "000011110010" => data <= X"204801D4";
         WHEN "000011110011" => data <= X"0418C3E2";
         WHEN "000011110100" => data <= X"042044E2";
         WHEN "000011110101" => data <= X"0000001A";
         WHEN "000011110110" => data <= X"0000801A";
         WHEN "000011110111" => data <= X"160000AB";
         WHEN "000011111000" => data <= X"200040AB";
         WHEN "000011111001" => data <= X"010080AB";
         WHEN "000011111010" => data <= X"0700C0AB";
         WHEN "000011111011" => data <= X"009094E5";
         WHEN "000011111100" => data <= X"0C000010";
         WHEN "000011111101" => data <= X"20002185";
         WHEN "000011111110" => data <= X"00000186";
         WHEN "000011111111" => data <= X"04004186";
         WHEN "000100000000" => data <= X"08008186";
         WHEN "000100000001" => data <= X"0C00C186";
         WHEN "000100000010" => data <= X"10000187";
         WHEN "000100000011" => data <= X"14004187";
         WHEN "000100000100" => data <= X"18008187";
         WHEN "000100000101" => data <= X"1C00C187";
         WHEN "000100000110" => data <= X"00480044";
         WHEN "000100000111" => data <= X"2400219C";
         WHEN "000100001000" => data <= X"02C11070";
         WHEN "000100001001" => data <= X"180020AA";
         WHEN "000100001010" => data <= X"008076E2";
         WHEN "000100001011" => data <= X"0000B386";
         WHEN "000100001100" => data <= X"0102B572";
         WHEN "000100001101" => data <= X"02891570";
         WHEN "000100001110" => data <= X"0100319E";
         WHEN "000100001111" => data <= X"00D031E4";
         WHEN "000100010000" => data <= X"FBFFFF13";
         WHEN "000100010001" => data <= X"0400739E";
         WHEN "000100010010" => data <= X"02F11C70";
         WHEN "000100010011" => data <= X"C1FFFF07";
         WHEN "000100010100" => data <= X"0800949E";
         WHEN "000100010101" => data <= X"E6FFFF03";
         WHEN "000100010110" => data <= X"2000109E";
         WHEN "000100010111" => data <= X"B4FF219C";
         WHEN "000100011000" => data <= X"00F08018";
         WHEN "000100011001" => data <= X"2000A0A8";
         WHEN "000100011010" => data <= X"0823849C";
         WHEN "000100011011" => data <= X"0C00619C";
         WHEN "000100011100" => data <= X"2C8001D4";
         WHEN "000100011101" => data <= X"309001D4";
         WHEN "000100011110" => data <= X"38B001D4";
         WHEN "000100011111" => data <= X"3CC001D4";
         WHEN "000100100000" => data <= X"40D001D4";
         WHEN "000100100001" => data <= X"44E001D4";
         WHEN "000100100010" => data <= X"484801D4";
         WHEN "000100100011" => data <= X"34A001D4";
         WHEN "000100100100" => data <= X"A7010004";
         WHEN "000100100101" => data <= X"00F0401A";
         WHEN "000100100110" => data <= X"00F0001A";
         WHEN "000100100111" => data <= X"B009529E";
         WHEN "000100101000" => data <= X"180B109E";
         WHEN "000100101001" => data <= X"00F0A018";
         WHEN "000100101010" => data <= X"311BA59C";
         WHEN "000100101011" => data <= X"049092E0";
         WHEN "000100101100" => data <= X"BC000004";
         WHEN "000100101101" => data <= X"048070E0";
         WHEN "000100101110" => data <= X"1F00201A";
         WHEN "000100101111" => data <= X"00F0C01A";
         WHEN "000100110000" => data <= X"0000601A";
         WHEN "000100110001" => data <= X"00FC31AA";
         WHEN "000100110010" => data <= X"0004001B";
         WHEN "000100110011" => data <= X"FFFF40AF";
         WHEN "000100110100" => data <= X"621BD69E";
         WHEN "000100110101" => data <= X"010080AB";
         WHEN "000100110110" => data <= X"0200A0AA";
         WHEN "000100110111" => data <= X"08A891E2";
         WHEN "000100111000" => data <= X"00C094E2";
         WHEN "000100111001" => data <= X"0000B486";
         WHEN "000100111010" => data <= X"00D015E4";
         WHEN "000100111011" => data <= X"1D000010";
         WHEN "000100111100" => data <= X"0100319E";
         WHEN "000100111101" => data <= X"0000201A";
         WHEN "000100111110" => data <= X"008813E4";
         WHEN "000100111111" => data <= X"10000010";
         WHEN "000101000000" => data <= X"04B0B6E0";
         WHEN "000101000001" => data <= X"00F0A018";
         WHEN "000101000010" => data <= X"541BA59C";
         WHEN "000101000011" => data <= X"049092E0";
         WHEN "000101000100" => data <= X"048070E0";
         WHEN "000101000101" => data <= X"30004186";
         WHEN "000101000110" => data <= X"2C000186";
         WHEN "000101000111" => data <= X"34008186";
         WHEN "000101001000" => data <= X"3800C186";
         WHEN "000101001001" => data <= X"3C000187";
         WHEN "000101001010" => data <= X"40004187";
         WHEN "000101001011" => data <= X"44008187";
         WHEN "000101001100" => data <= X"48002185";
         WHEN "000101001101" => data <= X"9B000000";
         WHEN "000101001110" => data <= X"4C00219C";
         WHEN "000101001111" => data <= X"049092E0";
         WHEN "000101010000" => data <= X"98000004";
         WHEN "000101010001" => data <= X"048070E0";
         WHEN "000101010010" => data <= X"90FFFF07";
         WHEN "000101010011" => data <= X"04A074E0";
         WHEN "000101010100" => data <= X"1F00201A";
         WHEN "000101010101" => data <= X"04E07CE2";
         WHEN "000101010110" => data <= X"00FC31AA";
         WHEN "000101010111" => data <= X"0100319E";
         WHEN "000101011000" => data <= X"2000A01A";
         WHEN "000101011001" => data <= X"00A831E4";
         WHEN "000101011010" => data <= X"DDFFFF13";
         WHEN "000101011011" => data <= X"0200A0AA";
         WHEN "000101011100" => data <= X"00F0A018";
         WHEN "000101011101" => data <= X"7E1BA59C";
         WHEN "000101011110" => data <= X"049092E0";
         WHEN "000101011111" => data <= X"89000004";
         WHEN "000101100000" => data <= X"048070E0";
         WHEN "000101100001" => data <= X"0C00819E";
         WHEN "000101100010" => data <= X"04A074E2";
         WHEN "000101100011" => data <= X"180020AA";
         WHEN "000101100100" => data <= X"2000E0AA";
         WHEN "000101100101" => data <= X"0000B386";
         WHEN "000101100110" => data <= X"0102B572";
         WHEN "000101100111" => data <= X"02891570";
         WHEN "000101101000" => data <= X"0100319E";
         WHEN "000101101001" => data <= X"00B831E4";
         WHEN "000101101010" => data <= X"FBFFFF13";
         WHEN "000101101011" => data <= X"0400739E";
         WHEN "000101101100" => data <= X"7F00201A";
         WHEN "000101101101" => data <= X"00F031AA";
         WHEN "000101101110" => data <= X"160060AA";
         WHEN "000101101111" => data <= X"02991170";
         WHEN "000101110000" => data <= X"010020AA";
         WHEN "000101110001" => data <= X"070060AA";
         WHEN "000101110010" => data <= X"02991170";
         WHEN "000101110011" => data <= X"61FFFF07";
         WHEN "000101110100" => data <= X"00000015";
         WHEN "000101110101" => data <= X"00F0A018";
         WHEN "000101110110" => data <= X"9F1BA59C";
         WHEN "000101110111" => data <= X"049092E0";
         WHEN "000101111000" => data <= X"70000004";
         WHEN "000101111001" => data <= X"048070E0";
         WHEN "000101111010" => data <= X"7F04201A";
         WHEN "000101111011" => data <= X"00F031AA";
         WHEN "000101111100" => data <= X"0000601A";
         WHEN "000101111101" => data <= X"080020AB";
         WHEN "000101111110" => data <= X"0000B186";
         WHEN "000101111111" => data <= X"0000F486";
         WHEN "000110000000" => data <= X"00A817E4";
         WHEN "000110000001" => data <= X"14000010";
         WHEN "000110000010" => data <= X"0400319E";
         WHEN "000110000011" => data <= X"00F0A018";
         WHEN "000110000100" => data <= X"08B801D4";
         WHEN "000110000101" => data <= X"04A801D4";
         WHEN "000110000110" => data <= X"009801D4";
         WHEN "000110000111" => data <= X"049092E0";
         WHEN "000110001000" => data <= X"048070E0";
         WHEN "000110001001" => data <= X"5F000004";
         WHEN "000110001010" => data <= X"C41BA59C";
         WHEN "000110001011" => data <= X"48002185";
         WHEN "000110001100" => data <= X"2C000186";
         WHEN "000110001101" => data <= X"30004186";
         WHEN "000110001110" => data <= X"34008186";
         WHEN "000110001111" => data <= X"3800C186";
         WHEN "000110010000" => data <= X"3C000187";
         WHEN "000110010001" => data <= X"40004187";
         WHEN "000110010010" => data <= X"44008187";
         WHEN "000110010011" => data <= X"00480044";
         WHEN "000110010100" => data <= X"4C00219C";
         WHEN "000110010101" => data <= X"0100739E";
         WHEN "000110010110" => data <= X"00C833E4";
         WHEN "000110010111" => data <= X"E7FFFF13";
         WHEN "000110011000" => data <= X"0400949E";
         WHEN "000110011001" => data <= X"00F0A018";
         WHEN "000110011010" => data <= X"A9FFFF03";
         WHEN "000110011011" => data <= X"E41BA59C";
         WHEN "000110011100" => data <= X"E8FF219C";
         WHEN "000110011101" => data <= X"008001D4";
         WHEN "000110011110" => data <= X"049001D4";
         WHEN "000110011111" => data <= X"08A001D4";
         WHEN "000110100000" => data <= X"0CB001D4";
         WHEN "000110100001" => data <= X"10C001D4";
         WHEN "000110100010" => data <= X"144801D4";
         WHEN "000110100011" => data <= X"041843E2";
         WHEN "000110100100" => data <= X"042084E2";
         WHEN "000110100101" => data <= X"1C0000AA";
         WHEN "000110100110" => data <= X"090000AB";
         WHEN "000110100111" => data <= X"FCFFC0AE";
         WHEN "000110101000" => data <= X"488074E0";
         WHEN "000110101001" => data <= X"0F0023A6";
         WHEN "000110101010" => data <= X"00C051E4";
         WHEN "000110101011" => data <= X"03000010";
         WHEN "000110101100" => data <= X"3700719C";
         WHEN "000110101101" => data <= X"3000719C";
         WHEN "000110101110" => data <= X"00900048";
         WHEN "000110101111" => data <= X"FCFF109E";
         WHEN "000110110000" => data <= X"00B030E4";
         WHEN "000110110001" => data <= X"F8FFFF13";
         WHEN "000110110010" => data <= X"488074E0";
         WHEN "000110110011" => data <= X"00000186";
         WHEN "000110110100" => data <= X"04004186";
         WHEN "000110110101" => data <= X"08008186";
         WHEN "000110110110" => data <= X"0C00C186";
         WHEN "000110110111" => data <= X"10000187";
         WHEN "000110111000" => data <= X"14002185";
         WHEN "000110111001" => data <= X"00480044";
         WHEN "000110111010" => data <= X"1800219C";
         WHEN "000110111011" => data <= X"E8FF219C";
         WHEN "000110111100" => data <= X"0C8001D4";
         WHEN "000110111101" => data <= X"109001D4";
         WHEN "000110111110" => data <= X"144801D4";
         WHEN "000110111111" => data <= X"041843E2";
         WHEN "000111000000" => data <= X"0000601A";
         WHEN "000111000001" => data <= X"0000001A";
         WHEN "000111000010" => data <= X"0A00A0AA";
         WHEN "000111000011" => data <= X"0AABE4E2";
         WHEN "000111000100" => data <= X"020020AA";
         WHEN "000111000101" => data <= X"088837E2";
         WHEN "000111000110" => data <= X"00B831E2";
         WHEN "000111000111" => data <= X"008831E2";
         WHEN "000111001000" => data <= X"028824E2";
         WHEN "000111001001" => data <= X"0200E19E";
         WHEN "000111001010" => data <= X"3000319E";
         WHEN "000111001011" => data <= X"0098F7E2";
         WHEN "000111001100" => data <= X"008817D8";
         WHEN "000111001101" => data <= X"0000201A";
         WHEN "000111001110" => data <= X"008813E4";
         WHEN "000111001111" => data <= X"04000010";
         WHEN "000111010000" => data <= X"008804E4";
         WHEN "000111010001" => data <= X"04000010";
         WHEN "000111010010" => data <= X"00000015";
         WHEN "000111010011" => data <= X"0100109E";
         WHEN "000111010100" => data <= X"FF0010A6";
         WHEN "000111010101" => data <= X"0100739E";
         WHEN "000111010110" => data <= X"00A833E4";
         WHEN "000111010111" => data <= X"ECFFFF13";
         WHEN "000111011000" => data <= X"0AAB84E0";
         WHEN "000111011001" => data <= X"0000201A";
         WHEN "000111011010" => data <= X"008830E4";
         WHEN "000111011011" => data <= X"07000010";
         WHEN "000111011100" => data <= X"FFFF109E";
         WHEN "000111011101" => data <= X"0C000186";
         WHEN "000111011110" => data <= X"10004186";
         WHEN "000111011111" => data <= X"14002185";
         WHEN "000111100000" => data <= X"00480044";
         WHEN "000111100001" => data <= X"1800219C";
         WHEN "000111100010" => data <= X"0200219E";
         WHEN "000111100011" => data <= X"008031E2";
         WHEN "000111100100" => data <= X"00900048";
         WHEN "000111100101" => data <= X"0000718C";
         WHEN "000111100110" => data <= X"F4FFFF03";
         WHEN "000111100111" => data <= X"0000201A";
         WHEN "000111101000" => data <= X"E0FF219C";
         WHEN "000111101001" => data <= X"008001D4";
         WHEN "000111101010" => data <= X"049001D4";
         WHEN "000111101011" => data <= X"08A001D4";
         WHEN "000111101100" => data <= X"0CB001D4";
         WHEN "000111101101" => data <= X"14D001D4";
         WHEN "000111101110" => data <= X"18E001D4";
         WHEN "000111101111" => data <= X"10C001D4";
         WHEN "000111110000" => data <= X"1C4801D4";
         WHEN "000111110001" => data <= X"041883E2";
         WHEN "000111110010" => data <= X"042004E2";
         WHEN "000111110011" => data <= X"042845E2";
         WHEN "000111110100" => data <= X"2000C19E";
         WHEN "000111110101" => data <= X"250040AB";
         WHEN "000111110110" => data <= X"630080AB";
         WHEN "000111110111" => data <= X"00007290";
         WHEN "000111111000" => data <= X"0000201A";
         WHEN "000111111001" => data <= X"008823E4";
         WHEN "000111111010" => data <= X"3B00000C";
         WHEN "000111111011" => data <= X"00D023E4";
         WHEN "000111111100" => data <= X"5A000010";
         WHEN "000111111101" => data <= X"FF0003A7";
         WHEN "000111111110" => data <= X"01003292";
         WHEN "000111111111" => data <= X"00E011E4";
         WHEN "001000000000" => data <= X"4D000010";
         WHEN "001000000001" => data <= X"00E051E5";
         WHEN "001000000010" => data <= X"1B000010";
         WHEN "001000000011" => data <= X"0000601A";
         WHEN "001000000100" => data <= X"009811E4";
         WHEN "001000000101" => data <= X"28000010";
         WHEN "001000000110" => data <= X"580060AA";
         WHEN "001000000111" => data <= X"009811E4";
         WHEN "001000001000" => data <= X"37000010";
         WHEN "001000001001" => data <= X"0400169F";
         WHEN "001000001010" => data <= X"00A00048";
         WHEN "001000001011" => data <= X"250060A8";
         WHEN "001000001100" => data <= X"0000201A";
         WHEN "001000001101" => data <= X"008810E4";
         WHEN "001000001110" => data <= X"04000010";
         WHEN "001000001111" => data <= X"00000015";
         WHEN "001000010000" => data <= X"00800048";
         WHEN "001000010001" => data <= X"250060A8";
         WHEN "001000010010" => data <= X"0100128F";
         WHEN "001000010011" => data <= X"00A00048";
         WHEN "001000010100" => data <= X"04C078E0";
         WHEN "001000010101" => data <= X"0000201A";
         WHEN "001000010110" => data <= X"008810E4";
         WHEN "001000010111" => data <= X"33000010";
         WHEN "001000011000" => data <= X"00000015";
         WHEN "001000011001" => data <= X"00800048";
         WHEN "001000011010" => data <= X"04C078E0";
         WHEN "001000011011" => data <= X"30000000";
         WHEN "001000011100" => data <= X"0100529E";
         WHEN "001000011101" => data <= X"640060AA";
         WHEN "001000011110" => data <= X"009811E4";
         WHEN "001000011111" => data <= X"EBFFFF0F";
         WHEN "001000100000" => data <= X"0400169F";
         WHEN "001000100001" => data <= X"04A074E0";
         WHEN "001000100010" => data <= X"0000D686";
         WHEN "001000100011" => data <= X"98FFFF07";
         WHEN "001000100100" => data <= X"04B096E0";
         WHEN "001000100101" => data <= X"0000201A";
         WHEN "001000100110" => data <= X"008810E4";
         WHEN "001000100111" => data <= X"22000010";
         WHEN "001000101000" => data <= X"04B096E0";
         WHEN "001000101001" => data <= X"92FFFF07";
         WHEN "001000101010" => data <= X"048070E0";
         WHEN "001000101011" => data <= X"1F000000";
         WHEN "001000101100" => data <= X"04C0D8E2";
         WHEN "001000101101" => data <= X"00A00048";
         WHEN "001000101110" => data <= X"04D07AE0";
         WHEN "001000101111" => data <= X"0000201A";
         WHEN "001000110000" => data <= X"008810E4";
         WHEN "001000110001" => data <= X"04000010";
         WHEN "001000110010" => data <= X"04D07AE0";
         WHEN "001000110011" => data <= X"00800048";
         WHEN "001000110100" => data <= X"00000015";
         WHEN "001000110101" => data <= X"00000186";
         WHEN "001000110110" => data <= X"04004186";
         WHEN "001000110111" => data <= X"08008186";
         WHEN "001000111000" => data <= X"0C00C186";
         WHEN "001000111001" => data <= X"10000187";
         WHEN "001000111010" => data <= X"14004187";
         WHEN "001000111011" => data <= X"18008187";
         WHEN "001000111100" => data <= X"1C002185";
         WHEN "001000111101" => data <= X"00480044";
         WHEN "001000111110" => data <= X"2000219C";
         WHEN "001000111111" => data <= X"04A074E0";
         WHEN "001001000000" => data <= X"0000D686";
         WHEN "001001000001" => data <= X"5BFFFF07";
         WHEN "001001000010" => data <= X"04B096E0";
         WHEN "001001000011" => data <= X"0000201A";
         WHEN "001001000100" => data <= X"008810E4";
         WHEN "001001000101" => data <= X"04000010";
         WHEN "001001000110" => data <= X"04B096E0";
         WHEN "001001000111" => data <= X"55FFFF07";
         WHEN "001001001000" => data <= X"048070E0";
         WHEN "001001001001" => data <= X"04C0D8E2";
         WHEN "001001001010" => data <= X"0100529E";
         WHEN "001001001011" => data <= X"ACFFFF03";
         WHEN "001001001100" => data <= X"0100529E";
         WHEN "001001001101" => data <= X"0300568E";
         WHEN "001001001110" => data <= X"00A00048";
         WHEN "001001001111" => data <= X"049072E0";
         WHEN "001001010000" => data <= X"0000201A";
         WHEN "001001010001" => data <= X"008810E4";
         WHEN "001001010010" => data <= X"E3FFFF13";
         WHEN "001001010011" => data <= X"049072E0";
         WHEN "001001010100" => data <= X"DFFFFF03";
         WHEN "001001010101" => data <= X"00000015";
         WHEN "001001010110" => data <= X"00A00048";
         WHEN "001001010111" => data <= X"04C078E0";
         WHEN "001001011000" => data <= X"0000201A";
         WHEN "001001011001" => data <= X"008810E4";
         WHEN "001001011010" => data <= X"F1FFFF13";
         WHEN "001001011011" => data <= X"00000015";
         WHEN "001001011100" => data <= X"00800048";
         WHEN "001001011101" => data <= X"04C078E0";
         WHEN "001001011110" => data <= X"99FFFF03";
         WHEN "001001011111" => data <= X"0100529E";
         WHEN "001001100000" => data <= X"0050201A";
         WHEN "001001100001" => data <= X"030071AA";
         WHEN "001001100010" => data <= X"83FFA0AE";
         WHEN "001001100011" => data <= X"00A813D8";
         WHEN "001001100100" => data <= X"1B00A0AA";
         WHEN "001001100101" => data <= X"00A811D8";
         WHEN "001001100110" => data <= X"010031AA";
         WHEN "001001100111" => data <= X"000011D8";
         WHEN "001001101000" => data <= X"030020AA";
         WHEN "001001101001" => data <= X"008813D8";
         WHEN "001001101010" => data <= X"00480044";
         WHEN "001001101011" => data <= X"00000015";
         WHEN "001001101100" => data <= X"0050601A";
         WHEN "001001101101" => data <= X"FF0063A4";
         WHEN "001001101110" => data <= X"0500B3AA";
         WHEN "001001101111" => data <= X"0000358E";
         WHEN "001001110000" => data <= X"400031A6";
         WHEN "001001110001" => data <= X"0000E01A";
         WHEN "001001110010" => data <= X"00B811E4";
         WHEN "001001110011" => data <= X"05000010";
         WHEN "001001110100" => data <= X"00000015";
         WHEN "001001110101" => data <= X"001813D8";
         WHEN "001001110110" => data <= X"00480044";
         WHEN "001001110111" => data <= X"00000015";
         WHEN "001001111000" => data <= X"00000015";
         WHEN "001001111001" => data <= X"F6FFFF03";
         WHEN "001001111010" => data <= X"00000015";
         WHEN "001001111011" => data <= X"0050601A";
         WHEN "001001111100" => data <= X"0500B3AA";
         WHEN "001001111101" => data <= X"0000358E";
         WHEN "001001111110" => data <= X"010031A6";
         WHEN "001001111111" => data <= X"0000E01A";
         WHEN "001010000000" => data <= X"00B811E4";
         WHEN "001010000001" => data <= X"FCFFFF13";
         WHEN "001010000010" => data <= X"00000015";
         WHEN "001010000011" => data <= X"0000738D";
         WHEN "001010000100" => data <= X"00480044";
         WHEN "001010000101" => data <= X"00000015";
         WHEN "001010000110" => data <= X"F0FF219C";
         WHEN "001010000111" => data <= X"FF0063A4";
         WHEN "001010001000" => data <= X"008001D4";
         WHEN "001010001001" => data <= X"D0FF039E";
         WHEN "001010001010" => data <= X"FF0030A6";
         WHEN "001010001011" => data <= X"090060AA";
         WHEN "001010001100" => data <= X"049001D4";
         WHEN "001010001101" => data <= X"08A001D4";
         WHEN "001010001110" => data <= X"009851E4";
         WHEN "001010001111" => data <= X"0800000C";
         WHEN "001010010000" => data <= X"0C4801D4";
         WHEN "001010010001" => data <= X"BFFF239E";
         WHEN "001010010010" => data <= X"FF0031A6";
         WHEN "001010010011" => data <= X"050060AA";
         WHEN "001010010100" => data <= X"009851E4";
         WHEN "001010010101" => data <= X"18000010";
         WHEN "001010010110" => data <= X"C9FF039E";
         WHEN "001010010111" => data <= X"090040AA";
         WHEN "001010011000" => data <= X"050080AA";
         WHEN "001010011001" => data <= X"E2FFFF07";
         WHEN "001010011010" => data <= X"00000015";
         WHEN "001010011011" => data <= X"FF006BA5";
         WHEN "001010011100" => data <= X"D0FF2B9E";
         WHEN "001010011101" => data <= X"FF0071A6";
         WHEN "001010011110" => data <= X"009053E4";
         WHEN "001010011111" => data <= X"04000010";
         WHEN "001010100000" => data <= X"0400A0AA";
         WHEN "001010100001" => data <= X"08A810E2";
         WHEN "001010100010" => data <= X"008011E2";
         WHEN "001010100011" => data <= X"BFFF2B9E";
         WHEN "001010100100" => data <= X"FF0031A6";
         WHEN "001010100101" => data <= X"00A051E4";
         WHEN "001010100110" => data <= X"10000010";
         WHEN "001010100111" => data <= X"9FFF2B9E";
         WHEN "001010101000" => data <= X"040020AA";
         WHEN "001010101001" => data <= X"088810E2";
         WHEN "001010101010" => data <= X"C9FF6B9D";
         WHEN "001010101011" => data <= X"EEFFFF03";
         WHEN "001010101100" => data <= X"00800BE2";
         WHEN "001010101101" => data <= X"9FFF239E";
         WHEN "001010101110" => data <= X"FF0031A6";
         WHEN "001010101111" => data <= X"009851E4";
         WHEN "001010110000" => data <= X"04000010";
         WHEN "001010110001" => data <= X"00000015";
         WHEN "001010110010" => data <= X"E5FFFF03";
         WHEN "001010110011" => data <= X"A9FF039E";
         WHEN "001010110100" => data <= X"E3FFFF03";
         WHEN "001010110101" => data <= X"0000001A";
         WHEN "001010110110" => data <= X"FF0031A6";
         WHEN "001010110111" => data <= X"00A051E4";
         WHEN "001010111000" => data <= X"05000010";
         WHEN "001010111001" => data <= X"040020AA";
         WHEN "001010111010" => data <= X"088810E2";
         WHEN "001010111011" => data <= X"F0FFFF03";
         WHEN "001010111100" => data <= X"A9FF6B9D";
         WHEN "001010111101" => data <= X"0090B3E4";
         WHEN "001010111110" => data <= X"DBFFFF13";
         WHEN "001010111111" => data <= X"048070E1";
         WHEN "001011000000" => data <= X"04004186";
         WHEN "001011000001" => data <= X"00000186";
         WHEN "001011000010" => data <= X"08008186";
         WHEN "001011000011" => data <= X"0C002185";
         WHEN "001011000100" => data <= X"00480044";
         WHEN "001011000101" => data <= X"1000219C";
         WHEN "001011000110" => data <= X"FF0063A4";
         WHEN "001011000111" => data <= X"020020AA";
         WHEN "001011001000" => data <= X"00191170";
         WHEN "001011001001" => data <= X"00480044";
         WHEN "001011001010" => data <= X"00000015";
         WHEN "001011001011" => data <= X"041863E1";
         WHEN "001011001100" => data <= X"0000201A";
         WHEN "001011001101" => data <= X"002831E4";
         WHEN "001011001110" => data <= X"04000010";
         WHEN "001011001111" => data <= X"008864E2";
         WHEN "001011010000" => data <= X"00480044";
         WHEN "001011010001" => data <= X"00000015";
         WHEN "001011010010" => data <= X"0000B392";
         WHEN "001011010011" => data <= X"00886BE2";
         WHEN "001011010100" => data <= X"00A813D8";
         WHEN "001011010101" => data <= X"F8FFFF03";
         WHEN "001011010110" => data <= X"0100319E";
         WHEN "001011010111" => data <= X"9CFF219C";
         WHEN "001011011000" => data <= X"00F08018";
         WHEN "001011011001" => data <= X"3C00A0A8";
         WHEN "001011011010" => data <= X"2823849C";
         WHEN "001011011011" => data <= X"4C8001D4";
         WHEN "001011011100" => data <= X"509001D4";
         WHEN "001011011101" => data <= X"54A001D4";
         WHEN "001011011110" => data <= X"58B001D4";
         WHEN "001011011111" => data <= X"5CC001D4";
         WHEN "001011100000" => data <= X"604801D4";
         WHEN "001011100001" => data <= X"EAFFFF07";
         WHEN "001011100010" => data <= X"1000619C";
         WHEN "001011100011" => data <= X"030020AA";
         WHEN "001011100100" => data <= X"00011170";
         WHEN "001011100101" => data <= X"FF0020AA";
         WHEN "001011100110" => data <= X"090000B6";
         WHEN "001011100111" => data <= X"0088B0E4";
         WHEN "001011101000" => data <= X"FEFFFF13";
         WHEN "001011101001" => data <= X"0F00D0A6";
         WHEN "001011101010" => data <= X"010020AA";
         WHEN "001011101011" => data <= X"008836E4";
         WHEN "001011101100" => data <= X"5C000010";
         WHEN "001011101101" => data <= X"00000015";
         WHEN "001011101110" => data <= X"00F0801A";
         WHEN "001011101111" => data <= X"B009949E";
         WHEN "001011110000" => data <= X"00F0401A";
         WHEN "001011110001" => data <= X"180B529E";
         WHEN "001011110010" => data <= X"00F0A018";
         WHEN "001011110011" => data <= X"04A094E0";
         WHEN "001011110100" => data <= X"F71BA59C";
         WHEN "001011110101" => data <= X"F3FEFF07";
         WHEN "001011110110" => data <= X"049072E0";
         WHEN "001011110111" => data <= X"00F0A018";
         WHEN "001011111000" => data <= X"04A094E0";
         WHEN "001011111001" => data <= X"261CA59C";
         WHEN "001011111010" => data <= X"EEFEFF07";
         WHEN "001011111011" => data <= X"049072E0";
         WHEN "001011111100" => data <= X"00F0A018";
         WHEN "001011111101" => data <= X"04A094E0";
         WHEN "001011111110" => data <= X"491CA59C";
         WHEN "001011111111" => data <= X"E9FEFF07";
         WHEN "001100000000" => data <= X"049072E0";
         WHEN "001100000001" => data <= X"040020AA";
         WHEN "001100000010" => data <= X"488830E2";
         WHEN "001100000011" => data <= X"0F0031A6";
         WHEN "001100000100" => data <= X"00F0A018";
         WHEN "001100000101" => data <= X"04A094E0";
         WHEN "001100000110" => data <= X"048801D4";
         WHEN "001100000111" => data <= X"7B1CA59C";
         WHEN "001100001000" => data <= X"049072E0";
         WHEN "001100001001" => data <= X"DFFEFF07";
         WHEN "001100001010" => data <= X"00B001D4";
         WHEN "001100001011" => data <= X"0C0020AA";
         WHEN "001100001100" => data <= X"488830E2";
         WHEN "001100001101" => data <= X"0F0031A6";
         WHEN "001100001110" => data <= X"0C8801D4";
         WHEN "001100001111" => data <= X"100020AA";
         WHEN "001100010000" => data <= X"488830E2";
         WHEN "001100010001" => data <= X"0F0031A6";
         WHEN "001100010010" => data <= X"088801D4";
         WHEN "001100010011" => data <= X"140020AA";
         WHEN "001100010100" => data <= X"488830E2";
         WHEN "001100010101" => data <= X"0F0031A6";
         WHEN "001100010110" => data <= X"048801D4";
         WHEN "001100010111" => data <= X"180020AA";
         WHEN "001100011000" => data <= X"488810E2";
         WHEN "001100011001" => data <= X"0F0010A6";
         WHEN "001100011010" => data <= X"00F0A018";
         WHEN "001100011011" => data <= X"008001D4";
         WHEN "001100011100" => data <= X"04A094E0";
         WHEN "001100011101" => data <= X"991CA59C";
         WHEN "001100011110" => data <= X"049072E0";
         WHEN "001100011111" => data <= X"C9FEFF07";
         WHEN "001100100000" => data <= X"00F0801A";
         WHEN "001100100001" => data <= X"1000019E";
         WHEN "001100100010" => data <= X"010000AB";
         WHEN "001100100011" => data <= X"B009949E";
         WHEN "001100100100" => data <= X"0000201A";
         WHEN "001100100101" => data <= X"0000B084";
         WHEN "001100100110" => data <= X"008825E4";
         WHEN "001100100111" => data <= X"23000010";
         WHEN "001100101000" => data <= X"00C016E4";
         WHEN "001100101001" => data <= X"00C036E4";
         WHEN "001100101010" => data <= X"1600000C";
         WHEN "001100101011" => data <= X"00000015";
         WHEN "001100101100" => data <= X"00F0A018";
         WHEN "001100101101" => data <= X"AA1CA59C";
         WHEN "001100101110" => data <= X"00008018";
         WHEN "001100101111" => data <= X"B9FEFF07";
         WHEN "001100110000" => data <= X"049072E0";
         WHEN "001100110001" => data <= X"025020B6";
         WHEN "001100110010" => data <= X"0000601A";
         WHEN "001100110011" => data <= X"009871E5";
         WHEN "001100110100" => data <= X"FDFFFF13";
         WHEN "001100110101" => data <= X"00000015";
         WHEN "001100110110" => data <= X"035000B6";
         WHEN "001100110111" => data <= X"00F0A018";
         WHEN "001100111000" => data <= X"008001D4";
         WHEN "001100111001" => data <= X"CC1CA59C";
         WHEN "001100111010" => data <= X"00008018";
         WHEN "001100111011" => data <= X"ADFEFF07";
         WHEN "001100111100" => data <= X"049072E0";
         WHEN "001100111101" => data <= X"00800044";
         WHEN "001100111110" => data <= X"00000015";
         WHEN "001100111111" => data <= X"00000015";
         WHEN "001101000000" => data <= X"4C000186";
         WHEN "001101000001" => data <= X"50004186";
         WHEN "001101000010" => data <= X"54008186";
         WHEN "001101000011" => data <= X"5800C186";
         WHEN "001101000100" => data <= X"5C000187";
         WHEN "001101000101" => data <= X"60002185";
         WHEN "001101000110" => data <= X"00480044";
         WHEN "001101000111" => data <= X"6400219C";
         WHEN "001101001000" => data <= X"A8FFFF03";
         WHEN "001101001001" => data <= X"0000801A";
         WHEN "001101001010" => data <= X"E2FFFF0F";
         WHEN "001101001011" => data <= X"0400109E";
         WHEN "001101001100" => data <= X"04A094E0";
         WHEN "001101001101" => data <= X"9BFEFF07";
         WHEN "001101001110" => data <= X"049072E0";
         WHEN "001101001111" => data <= X"D6FFFF03";
         WHEN "001101010000" => data <= X"0000201A";
         WHEN "001101010001" => data <= X"ADDE201A";
         WHEN "001101010010" => data <= X"001371AA";
         WHEN "001101010011" => data <= X"009803E4";
         WHEN "001101010100" => data <= X"13000010";
         WHEN "001101010101" => data <= X"FFFF601A";
         WHEN "001101010110" => data <= X"039863E0";
         WHEN "001101010111" => data <= X"008823E4";
         WHEN "001101011000" => data <= X"10000010";
         WHEN "001101011001" => data <= X"FFFF60AD";
         WHEN "001101011010" => data <= X"00F0A018";
         WHEN "001101011011" => data <= X"00F08018";
         WHEN "001101011100" => data <= X"00F06018";
         WHEN "001101011101" => data <= X"FCFF219C";
         WHEN "001101011110" => data <= X"EB1CA59C";
         WHEN "001101011111" => data <= X"B009849C";
         WHEN "001101100000" => data <= X"004801D4";
         WHEN "001101100001" => data <= X"87FEFF07";
         WHEN "001101100010" => data <= X"180B639C";
         WHEN "001101100011" => data <= X"FFFF60AD";
         WHEN "001101100100" => data <= X"00002185";
         WHEN "001101100101" => data <= X"00480044";
         WHEN "001101100110" => data <= X"0400219C";
         WHEN "001101100111" => data <= X"00006019";
         WHEN "001101101000" => data <= X"00480044";
         WHEN "001101101001" => data <= X"00000015";
         WHEN "001101101010" => data <= X"A4FC219C";
         WHEN "001101101011" => data <= X"307301D4";
         WHEN "001101101100" => data <= X"348301D4";
         WHEN "001101101101" => data <= X"389301D4";
         WHEN "001101101110" => data <= X"3CA301D4";
         WHEN "001101101111" => data <= X"40B301D4";
         WHEN "001101110000" => data <= X"44C301D4";
         WHEN "001101110001" => data <= X"48D301D4";
         WHEN "001101110010" => data <= X"4CE301D4";
         WHEN "001101110011" => data <= X"50F301D4";
         WHEN "001101110100" => data <= X"541301D4";
         WHEN "001101110101" => data <= X"584B01D4";
         WHEN "001101110110" => data <= X"00C0201A";
         WHEN "001101110111" => data <= X"068800C0";
         WHEN "001101111000" => data <= X"110020B6";
         WHEN "001101111001" => data <= X"2C8801D4";
         WHEN "001101111010" => data <= X"2C002186";
         WHEN "001101111011" => data <= X"100031AA";
         WHEN "001101111100" => data <= X"2C8801D4";
         WHEN "001101111101" => data <= X"2C002186";
         WHEN "001101111110" => data <= X"118800C0";
         WHEN "001101111111" => data <= X"E1FEFF07";
         WHEN "001110000000" => data <= X"7F00C01B";
         WHEN "001110000001" => data <= X"56FFFF07";
         WHEN "001110000010" => data <= X"010040AA";
         WHEN "001110000011" => data <= X"00F0201A";
         WHEN "001110000100" => data <= X"004031AA";
         WHEN "001110000101" => data <= X"108801D4";
         WHEN "001110000110" => data <= X"3F00201A";
         WHEN "001110000111" => data <= X"FFFF31AA";
         WHEN "001110001000" => data <= X"FCFFDEAB";
         WHEN "001110001001" => data <= X"0000C019";
         WHEN "001110001010" => data <= X"0000001B";
         WHEN "001110001011" => data <= X"049052E0";
         WHEN "001110001100" => data <= X"0000001A";
         WHEN "001110001101" => data <= X"1C8801D4";
         WHEN "001110001110" => data <= X"270080AB";
         WHEN "001110001111" => data <= X"ECFEFF07";
         WHEN "001110010000" => data <= X"00000015";
         WHEN "001110010001" => data <= X"FF004BA7";
         WHEN "001110010010" => data <= X"00E01AE4";
         WHEN "001110010011" => data <= X"AF020010";
         WHEN "001110010100" => data <= X"00E05AE4";
         WHEN "001110010101" => data <= X"4A000010";
         WHEN "001110010110" => data <= X"240020AA";
         WHEN "001110010111" => data <= X"00881AE4";
         WHEN "001110011000" => data <= X"A2000010";
         WHEN "001110011001" => data <= X"00885AE4";
         WHEN "001110011010" => data <= X"13000010";
         WHEN "001110011011" => data <= X"230020AA";
         WHEN "001110011100" => data <= X"00881AE4";
         WHEN "001110011101" => data <= X"93000010";
         WHEN "001110011110" => data <= X"F6FF7A9E";
         WHEN "001110011111" => data <= X"FF0073A6";
         WHEN "001110100000" => data <= X"160020AA";
         WHEN "001110100001" => data <= X"008853E4";
         WHEN "001110100010" => data <= X"09000010";
         WHEN "001110100011" => data <= X"BFFF201A";
         WHEN "001110100100" => data <= X"F6FF31AA";
         WHEN "001110100101" => data <= X"889831E2";
         WHEN "001110100110" => data <= X"010031A6";
         WHEN "001110100111" => data <= X"0000601A";
         WHEN "001110101000" => data <= X"009831E4";
         WHEN "001110101001" => data <= X"E6FFFF0F";
         WHEN "001110101010" => data <= X"00000015";
         WHEN "001110101011" => data <= X"46000000";
         WHEN "001110101100" => data <= X"00006019";
         WHEN "001110101101" => data <= X"260020AA";
         WHEN "001110101110" => data <= X"00881AE4";
         WHEN "001110101111" => data <= X"FCFFFF0F";
         WHEN "001110110000" => data <= X"250040AB";
         WHEN "001110110001" => data <= X"CAFEFF07";
         WHEN "001110110010" => data <= X"0000801B";
         WHEN "001110110011" => data <= X"00F0A018";
         WHEN "001110110100" => data <= X"00F06018";
         WHEN "001110110101" => data <= X"FF006BA5";
         WHEN "001110110110" => data <= X"4D1DA59C";
         WHEN "001110110111" => data <= X"00008018";
         WHEN "001110111000" => data <= X"180B639C";
         WHEN "001110111001" => data <= X"2FFEFF07";
         WHEN "001110111010" => data <= X"0C5801D4";
         WHEN "001110111011" => data <= X"200040AB";
         WHEN "001110111100" => data <= X"0C006185";
         WHEN "001110111101" => data <= X"00D00BE4";
         WHEN "001110111110" => data <= X"1D000010";
         WHEN "001110111111" => data <= X"00E03CE2";
         WHEN "001111000000" => data <= X"00E031E2";
         WHEN "001111000001" => data <= X"3000619E";
         WHEN "001111000010" => data <= X"0088F3E2";
         WHEN "001111000011" => data <= X"0000A01A";
         WHEN "001111000100" => data <= X"0100B59E";
         WHEN "001111000101" => data <= X"005817D8";
         WHEN "001111000110" => data <= X"188801D4";
         WHEN "001111000111" => data <= X"14A801D4";
         WHEN "001111001000" => data <= X"B3FEFF07";
         WHEN "001111001001" => data <= X"0CB801D4";
         WHEN "001111001010" => data <= X"FF006BA5";
         WHEN "001111001011" => data <= X"00D02BE4";
         WHEN "001111001100" => data <= X"0C00E186";
         WHEN "001111001101" => data <= X"1400A186";
         WHEN "001111001110" => data <= X"0100F79E";
         WHEN "001111001111" => data <= X"F5FFFF13";
         WHEN "001111010000" => data <= X"18002186";
         WHEN "001111010001" => data <= X"1003319E";
         WHEN "001111010010" => data <= X"2000619E";
         WHEN "001111010011" => data <= X"009831E2";
         WHEN "001111010100" => data <= X"00A831E2";
         WHEN "001111010101" => data <= X"0005F1DB";
         WHEN "001111010110" => data <= X"01009C9F";
         WHEN "001111010111" => data <= X"FF0020AA";
         WHEN "001111011000" => data <= X"0088BCE5";
         WHEN "001111011001" => data <= X"B5FFFF0F";
         WHEN "001111011010" => data <= X"00000015";
         WHEN "001111011011" => data <= X"A0FEFF07";
         WHEN "001111011100" => data <= X"00000015";
         WHEN "001111011101" => data <= X"E0FFFF03";
         WHEN "001111011110" => data <= X"FF006BA5";
         WHEN "001111011111" => data <= X"2D0020AA";
         WHEN "001111100000" => data <= X"00881AE4";
         WHEN "001111100001" => data <= X"0B000010";
         WHEN "001111100010" => data <= X"00885AE4";
         WHEN "001111100011" => data <= X"33000010";
         WHEN "001111100100" => data <= X"3D0020AA";
         WHEN "001111100101" => data <= X"2A0020AA";
         WHEN "001111100110" => data <= X"00881AE4";
         WHEN "001111100111" => data <= X"7F000010";
         WHEN "001111101000" => data <= X"2B0020AA";
         WHEN "001111101001" => data <= X"00881AE4";
         WHEN "001111101010" => data <= X"0700000C";
         WHEN "001111101011" => data <= X"00006019";
         WHEN "001111101100" => data <= X"8FFEFF07";
         WHEN "001111101101" => data <= X"00000015";
         WHEN "001111101110" => data <= X"180020AA";
         WHEN "001111101111" => data <= X"08886BE1";
         WHEN "001111110000" => data <= X"88886BE1";
         WHEN "001111110001" => data <= X"180020AA";
         WHEN "001111110010" => data <= X"08885AE3";
         WHEN "001111110011" => data <= X"88885AE3";
         WHEN "001111110100" => data <= X"FFFF80AF";
         WHEN "001111110101" => data <= X"0000201A";
         WHEN "001111110110" => data <= X"FF00A0AA";
         WHEN "001111110111" => data <= X"008871E2";
         WHEN "001111111000" => data <= X"008873E2";
         WHEN "001111111001" => data <= X"2000E19E";
         WHEN "001111111010" => data <= X"1003739E";
         WHEN "001111111011" => data <= X"00B873E2";
         WHEN "001111111100" => data <= X"00FDF392";
         WHEN "001111111101" => data <= X"00D037E4";
         WHEN "001111111110" => data <= X"08000010";
         WHEN "001111111111" => data <= X"00000015";
         WHEN "010000000000" => data <= X"01FD7392";
         WHEN "010000000001" => data <= X"005813E4";
         WHEN "010000000010" => data <= X"0400000C";
         WHEN "010000000011" => data <= X"00000015";
         WHEN "010000000100" => data <= X"048891E3";
         WHEN "010000000101" => data <= X"000120AA";
         WHEN "010000000110" => data <= X"0100319E";
         WHEN "010000000111" => data <= X"00A8B1E5";
         WHEN "010000001000" => data <= X"F0FFFF13";
         WHEN "010000001001" => data <= X"008871E2";
         WHEN "010000001010" => data <= X"0000201A";
         WHEN "010000001011" => data <= X"00887CE5";
         WHEN "010000001100" => data <= X"4302000C";
         WHEN "010000001101" => data <= X"00F0A018";
         WHEN "010000001110" => data <= X"00F0201A";
         WHEN "010000001111" => data <= X"D820519F";
         WHEN "010000010000" => data <= X"0000201A";
         WHEN "010000010001" => data <= X"008832E4";
         WHEN "010000010010" => data <= X"40020010";
         WHEN "010000010011" => data <= X"00880EE4";
         WHEN "010000010100" => data <= X"7AFFFF03";
         WHEN "010000010101" => data <= X"010040AA";
         WHEN "010000010110" => data <= X"00881AE4";
         WHEN "010000010111" => data <= X"D5FFFF13";
         WHEN "010000011000" => data <= X"400020AA";
         WHEN "010000011001" => data <= X"00881AE4";
         WHEN "010000011010" => data <= X"D7FFFF0F";
         WHEN "010000011011" => data <= X"00006019";
         WHEN "010000011100" => data <= X"6AFEFF07";
         WHEN "010000011101" => data <= X"200060A8";
         WHEN "010000011110" => data <= X"020020AA";
         WHEN "010000011111" => data <= X"00F0A018";
         WHEN "010000100000" => data <= X"00F06018";
         WHEN "010000100001" => data <= X"48888BE2";
         WHEN "010000100010" => data <= X"005801D4";
         WHEN "010000100011" => data <= X"1C002186";
         WHEN "010000100100" => data <= X"611DA59C";
         WHEN "010000100101" => data <= X"00008018";
         WHEN "010000100110" => data <= X"180B639C";
         WHEN "010000100111" => data <= X"038894E2";
         WHEN "010000101000" => data <= X"C0FDFF07";
         WHEN "010000101001" => data <= X"0458CBE2";
         WHEN "010000101010" => data <= X"0000201A";
         WHEN "010000101011" => data <= X"008814E4";
         WHEN "010000101100" => data <= X"62FFFF0F";
         WHEN "010000101101" => data <= X"0000C019";
         WHEN "010000101110" => data <= X"60FFFF03";
         WHEN "010000101111" => data <= X"0000001B";
         WHEN "010000110000" => data <= X"00F0A018";
         WHEN "010000110001" => data <= X"3D1DA59C";
         WHEN "010000110010" => data <= X"00F08018";
         WHEN "010000110011" => data <= X"B009849C";
         WHEN "010000110100" => data <= X"00F06018";
         WHEN "010000110101" => data <= X"180B639C";
         WHEN "010000110110" => data <= X"B2FDFF07";
         WHEN "010000110111" => data <= X"270080AB";
         WHEN "010000111000" => data <= X"57FFFF03";
         WHEN "010000111001" => data <= X"00000015";
         WHEN "010000111010" => data <= X"00007084";
         WHEN "010000111011" => data <= X"16FFFF07";
         WHEN "010000111100" => data <= X"00000015";
         WHEN "010000111101" => data <= X"0000201A";
         WHEN "010000111110" => data <= X"00880BE4";
         WHEN "010000111111" => data <= X"05000010";
         WHEN "010001000000" => data <= X"10002186";
         WHEN "010001000001" => data <= X"00F0A018";
         WHEN "010001000010" => data <= X"F0FFFF03";
         WHEN "010001000011" => data <= X"7F1DA59C";
         WHEN "010001000100" => data <= X"008830E4";
         WHEN "010001000101" => data <= X"05000010";
         WHEN "010001000110" => data <= X"010020AA";
         WHEN "010001000111" => data <= X"0F8880C3";
         WHEN "010001001000" => data <= X"47FFFF03";
         WHEN "010001001001" => data <= X"270080AB";
         WHEN "010001001010" => data <= X"110020B6";
         WHEN "010001001011" => data <= X"FFBF60AE";
         WHEN "010001001100" => data <= X"2C8801D4";
         WHEN "010001001101" => data <= X"2C002186";
         WHEN "010001001110" => data <= X"039831E2";
         WHEN "010001001111" => data <= X"2C8801D4";
         WHEN "010001010000" => data <= X"20F040C1";
         WHEN "010001010001" => data <= X"2C002186";
         WHEN "010001010010" => data <= X"118800C0";
         WHEN "010001010011" => data <= X"E7BF60AE";
         WHEN "010001010100" => data <= X"2C002186";
         WHEN "010001010101" => data <= X"039831E2";
         WHEN "010001010110" => data <= X"2C8801D4";
         WHEN "010001010111" => data <= X"0D0040AB";
         WHEN "010001011000" => data <= X"00E05AB7";
         WHEN "010001011001" => data <= X"00F0A018";
         WHEN "010001011010" => data <= X"00F08018";
         WHEN "010001011011" => data <= X"00F06018";
         WHEN "010001011100" => data <= X"9A1DA59C";
         WHEN "010001011101" => data <= X"B009849C";
         WHEN "010001011110" => data <= X"8AFDFF07";
         WHEN "010001011111" => data <= X"180B639C";
         WHEN "010001100000" => data <= X"04D050E3";
         WHEN "010001100001" => data <= X"2C002186";
         WHEN "010001100010" => data <= X"00D00044";
         WHEN "010001100011" => data <= X"118800C0";
         WHEN "010001100100" => data <= X"2BFFFF03";
         WHEN "010001100101" => data <= X"270080AB";
         WHEN "010001100110" => data <= X"15FEFF07";
         WHEN "010001100111" => data <= X"00000015";
         WHEN "010001101000" => data <= X"FF006BA5";
         WHEN "010001101001" => data <= X"700020AA";
         WHEN "010001101010" => data <= X"00880BE4";
         WHEN "010001101011" => data <= X"CE000010";
         WHEN "010001101100" => data <= X"00884BE4";
         WHEN "010001101101" => data <= X"7A000010";
         WHEN "010001101110" => data <= X"680020AA";
         WHEN "010001101111" => data <= X"00880BE4";
         WHEN "010001110000" => data <= X"9D000010";
         WHEN "010001110001" => data <= X"00884BE4";
         WHEN "010001110010" => data <= X"15000010";
         WHEN "010001110011" => data <= X"650020AA";
         WHEN "010001110100" => data <= X"00880BE4";
         WHEN "010001110101" => data <= X"96010010";
         WHEN "010001110110" => data <= X"660020AA";
         WHEN "010001110111" => data <= X"00880BE4";
         WHEN "010001111000" => data <= X"3C010010";
         WHEN "010001111001" => data <= X"630020AA";
         WHEN "010001111010" => data <= X"00880BE4";
         WHEN "010001111011" => data <= X"13FFFF0F";
         WHEN "010001111100" => data <= X"00F0201A";
         WHEN "010001111101" => data <= X"004031AA";
         WHEN "010001111110" => data <= X"008810E4";
         WHEN "010001111111" => data <= X"05000010";
         WHEN "010010000000" => data <= X"0004201A";
         WHEN "010010000001" => data <= X"008830E4";
         WHEN "010010000010" => data <= X"FB000010";
         WHEN "010010000011" => data <= X"00000015";
         WHEN "010010000100" => data <= X"00F0A018";
         WHEN "010010000101" => data <= X"ADFFFF03";
         WHEN "010010000110" => data <= X"681EA59C";
         WHEN "010010000111" => data <= X"690020AA";
         WHEN "010010001000" => data <= X"00880BE4";
         WHEN "010010001001" => data <= X"B9000010";
         WHEN "010010001010" => data <= X"6D0020AA";
         WHEN "010010001011" => data <= X"00880BE4";
         WHEN "010010001100" => data <= X"02FFFF0F";
         WHEN "010010001101" => data <= X"00F0401B";
         WHEN "010010001110" => data <= X"00F0001B";
         WHEN "010010001111" => data <= X"180B389E";
         WHEN "010010010000" => data <= X"B0095A9F";
         WHEN "010010010001" => data <= X"00F0A018";
         WHEN "010010010010" => data <= X"048871E0";
         WHEN "010010010011" => data <= X"AD1FA59C";
         WHEN "010010010100" => data <= X"04D09AE0";
         WHEN "010010010101" => data <= X"53FDFF07";
         WHEN "010010010110" => data <= X"0C8801D4";
         WHEN "010010010111" => data <= X"00F0201A";
         WHEN "010010011000" => data <= X"CF1F319E";
         WHEN "010010011001" => data <= X"148801D4";
         WHEN "010010011010" => data <= X"00F0201A";
         WHEN "010010011011" => data <= X"E91F319E";
         WHEN "010010011100" => data <= X"0000001B";
         WHEN "010010011101" => data <= X"188801D4";
         WHEN "010010011110" => data <= X"04D09AE0";
         WHEN "010010011111" => data <= X"1400A184";
         WHEN "010010100000" => data <= X"48FDFF07";
         WHEN "010010100001" => data <= X"0C006184";
         WHEN "010010100010" => data <= X"0000201A";
         WHEN "010010100011" => data <= X"0002601A";
         WHEN "010010100100" => data <= X"0200A0AA";
         WHEN "010010100101" => data <= X"00A818E4";
         WHEN "010010100110" => data <= X"03000010";
         WHEN "010010100111" => data <= X"00000015";
         WHEN "010010101000" => data <= X"0100F172";
         WHEN "010010101001" => data <= X"008811D4";
         WHEN "010010101010" => data <= X"0400319E";
         WHEN "010010101011" => data <= X"009831E4";
         WHEN "010010101100" => data <= X"F9FFFF13";
         WHEN "010010101101" => data <= X"0200A0AA";
         WHEN "010010101110" => data <= X"00F0A018";
         WHEN "010010101111" => data <= X"DB1FA59C";
         WHEN "010010110000" => data <= X"04D09AE0";
         WHEN "010010110001" => data <= X"37FDFF07";
         WHEN "010010110010" => data <= X"0C006184";
         WHEN "010010110011" => data <= X"0000201A";
         WHEN "010010110100" => data <= X"0000801B";
         WHEN "010010110101" => data <= X"1D0020AB";
         WHEN "010010110110" => data <= X"0002E01A";
         WHEN "010010110111" => data <= X"020060AA";
         WHEN "010010111000" => data <= X"009818E4";
         WHEN "010010111001" => data <= X"03000010";
         WHEN "010010111010" => data <= X"00000015";
         WHEN "010010111011" => data <= X"01007173";
         WHEN "010010111100" => data <= X"00007187";
         WHEN "010010111101" => data <= X"00881BE4";
         WHEN "010010111110" => data <= X"13000010";
         WHEN "010010111111" => data <= X"00C85CE4";
         WHEN "010011000000" => data <= X"10000010";
         WHEN "010011000001" => data <= X"00000015";
         WHEN "010011000010" => data <= X"00007187";
         WHEN "010011000011" => data <= X"04D09AE0";
         WHEN "010011000100" => data <= X"088801D4";
         WHEN "010011000101" => data <= X"008801D4";
         WHEN "010011000110" => data <= X"04D801D4";
         WHEN "010011000111" => data <= X"28C801D4";
         WHEN "010011001000" => data <= X"24B801D4";
         WHEN "010011001001" => data <= X"208801D4";
         WHEN "010011001010" => data <= X"1800A184";
         WHEN "010011001011" => data <= X"1DFDFF07";
         WHEN "010011001100" => data <= X"0C006184";
         WHEN "010011001101" => data <= X"28002187";
         WHEN "010011001110" => data <= X"2400E186";
         WHEN "010011001111" => data <= X"20002186";
         WHEN "010011010000" => data <= X"01009C9F";
         WHEN "010011010001" => data <= X"0400319E";
         WHEN "010011010010" => data <= X"00B831E4";
         WHEN "010011010011" => data <= X"E5FFFF13";
         WHEN "010011010100" => data <= X"020060AA";
         WHEN "010011010101" => data <= X"0000201A";
         WHEN "010011010110" => data <= X"00881CE4";
         WHEN "010011010111" => data <= X"60010010";
         WHEN "010011011000" => data <= X"030020AA";
         WHEN "010011011001" => data <= X"00F0A018";
         WHEN "010011011010" => data <= X"00E001D4";
         WHEN "010011011011" => data <= X"0520A59C";
         WHEN "010011011100" => data <= X"04D09AE0";
         WHEN "010011011101" => data <= X"0BFDFF07";
         WHEN "010011011110" => data <= X"0C006184";
         WHEN "010011011111" => data <= X"00F0A018";
         WHEN "010011100000" => data <= X"00E001D4";
         WHEN "010011100001" => data <= X"1E20A59C";
         WHEN "010011100010" => data <= X"04D09AE0";
         WHEN "010011100011" => data <= X"05FDFF07";
         WHEN "010011100100" => data <= X"0C006184";
         WHEN "010011100101" => data <= X"A9FEFF03";
         WHEN "010011100110" => data <= X"0000001B";
         WHEN "010011100111" => data <= X"730020AA";
         WHEN "010011101000" => data <= X"00880BE4";
         WHEN "010011101001" => data <= X"2E000010";
         WHEN "010011101010" => data <= X"00884BE4";
         WHEN "010011101011" => data <= X"14000010";
         WHEN "010011101100" => data <= X"740020AA";
         WHEN "010011101101" => data <= X"710020AA";
         WHEN "010011101110" => data <= X"00880BE4";
         WHEN "010011101111" => data <= X"2C00000C";
         WHEN "010011110000" => data <= X"0004401B";
         WHEN "010011110001" => data <= X"7F00401B";
         WHEN "010011110010" => data <= X"FCFF5AAB";
         WHEN "010011110011" => data <= X"00F08018";
         WHEN "010011110100" => data <= X"00F06018";
         WHEN "010011110101" => data <= X"00D03EE4";
         WHEN "010011110110" => data <= X"B009849C";
         WHEN "010011110111" => data <= X"46010010";
         WHEN "010011111000" => data <= X"180B639C";
         WHEN "010011111001" => data <= X"00F0A018";
         WHEN "010011111010" => data <= X"3920A59C";
         WHEN "010011111011" => data <= X"EDFCFF07";
         WHEN "010011111100" => data <= X"00C0C01B";
         WHEN "010011111101" => data <= X"91FEFF03";
         WHEN "010011111110" => data <= X"FC1FDEAB";
         WHEN "010011111111" => data <= X"00880BE4";
         WHEN "010100000000" => data <= X"5E000010";
         WHEN "010100000001" => data <= X"760020AA";
         WHEN "010100000010" => data <= X"00880BE4";
         WHEN "010100000011" => data <= X"8BFEFF0F";
         WHEN "010100000100" => data <= X"00F0A018";
         WHEN "010100000101" => data <= X"00F08018";
         WHEN "010100000110" => data <= X"00F06018";
         WHEN "010100000111" => data <= X"E01DA59C";
         WHEN "010100001000" => data <= X"B009849C";
         WHEN "010100001001" => data <= X"DFFCFF07";
         WHEN "010100001010" => data <= X"180B639C";
         WHEN "010100001011" => data <= X"83FEFF03";
         WHEN "010100001100" => data <= X"00004018";
         WHEN "010100001101" => data <= X"00F0A018";
         WHEN "010100001110" => data <= X"00F06018";
         WHEN "010100001111" => data <= X"AA1FA59C";
         WHEN "010100010000" => data <= X"00008018";
         WHEN "010100010001" => data <= X"D7FCFF07";
         WHEN "010100010010" => data <= X"B009639C";
         WHEN "010100010011" => data <= X"C4FDFF07";
         WHEN "010100010100" => data <= X"270080AB";
         WHEN "010100010101" => data <= X"7AFEFF03";
         WHEN "010100010110" => data <= X"00000015";
         WHEN "010100010111" => data <= X"00FCFF07";
         WHEN "010100011000" => data <= X"270080AB";
         WHEN "010100011001" => data <= X"76FEFF03";
         WHEN "010100011010" => data <= X"00000015";
         WHEN "010100011011" => data <= X"00007A84";
         WHEN "010100011100" => data <= X"35FEFF07";
         WHEN "010100011101" => data <= X"00000015";
         WHEN "010100011110" => data <= X"0000201A";
         WHEN "010100011111" => data <= X"00880BE4";
         WHEN "010100100000" => data <= X"04000010";
         WHEN "010100100001" => data <= X"00F0A018";
         WHEN "010100100010" => data <= X"10FFFF03";
         WHEN "010100100011" => data <= X"AF1DA59C";
         WHEN "010100100100" => data <= X"04003AAA";
         WHEN "010100100101" => data <= X"00007186";
         WHEN "010100100110" => data <= X"020020AA";
         WHEN "010100100111" => data <= X"088873E2";
         WHEN "010100101000" => data <= X"0000201A";
         WHEN "010100101001" => data <= X"008833E4";
         WHEN "010100101010" => data <= X"0A000010";
         WHEN "010100101011" => data <= X"0088BAE2";
         WHEN "010100101100" => data <= X"110020B6";
         WHEN "010100101101" => data <= X"FFBF60AE";
         WHEN "010100101110" => data <= X"2C8801D4";
         WHEN "010100101111" => data <= X"2C002186";
         WHEN "010100110000" => data <= X"039831E2";
         WHEN "010100110001" => data <= X"2C8801D4";
         WHEN "010100110010" => data <= X"1FFFFF03";
         WHEN "010100110011" => data <= X"00000015";
         WHEN "010100110100" => data <= X"0000B586";
         WHEN "010100110101" => data <= X"0400319E";
         WHEN "010100110110" => data <= X"FCAFF1D7";
         WHEN "010100110111" => data <= X"F3FFFF03";
         WHEN "010100111000" => data <= X"008833E4";
         WHEN "010100111001" => data <= X"00F0A018";
         WHEN "010100111010" => data <= X"00F08018";
         WHEN "010100111011" => data <= X"00F06018";
         WHEN "010100111100" => data <= X"CC1DA59C";
         WHEN "010100111101" => data <= X"B009849C";
         WHEN "010100111110" => data <= X"AAFCFF07";
         WHEN "010100111111" => data <= X"180B639C";
         WHEN "010101000000" => data <= X"4EFEFF03";
         WHEN "010101000001" => data <= X"010040A8";
         WHEN "010101000010" => data <= X"00007084";
         WHEN "010101000011" => data <= X"0EFEFF07";
         WHEN "010101000100" => data <= X"00000015";
         WHEN "010101000101" => data <= X"0000201A";
         WHEN "010101000110" => data <= X"00880BE4";
         WHEN "010101000111" => data <= X"00F08018";
         WHEN "010101001000" => data <= X"00F06018";
         WHEN "010101001001" => data <= X"04003086";
         WHEN "010101001010" => data <= X"B009849C";
         WHEN "010101001011" => data <= X"0A000010";
         WHEN "010101001100" => data <= X"180B639C";
         WHEN "010101001101" => data <= X"00F0A018";
         WHEN "010101001110" => data <= X"048801D4";
         WHEN "010101001111" => data <= X"000001D4";
         WHEN "010101010000" => data <= X"F51DA59C";
         WHEN "010101010001" => data <= X"97FCFF07";
         WHEN "010101010010" => data <= X"270080AB";
         WHEN "010101010011" => data <= X"3CFEFF03";
         WHEN "010101010100" => data <= X"00000015";
         WHEN "010101010101" => data <= X"020060AA";
         WHEN "010101010110" => data <= X"089831E2";
         WHEN "010101010111" => data <= X"048031E2";
         WHEN "010101011000" => data <= X"FFFF319E";
         WHEN "010101011001" => data <= X"00F0A018";
         WHEN "010101011010" => data <= X"048801D4";
         WHEN "010101011011" => data <= X"008001D4";
         WHEN "010101011100" => data <= X"F5FFFF03";
         WHEN "010101011101" => data <= X"091EA59C";
         WHEN "010101011110" => data <= X"0000201A";
         WHEN "010101011111" => data <= X"00F08018";
         WHEN "010101100000" => data <= X"00F06018";
         WHEN "010101100001" => data <= X"008830E4";
         WHEN "010101100010" => data <= X"B009849C";
         WHEN "010101100011" => data <= X"09000010";
         WHEN "010101100100" => data <= X"180B639C";
         WHEN "010101100101" => data <= X"00F0A018";
         WHEN "010101100110" => data <= X"2B1EA59C";
         WHEN "010101100111" => data <= X"81FCFF07";
         WHEN "010101101000" => data <= X"00F0001A";
         WHEN "010101101001" => data <= X"0000001B";
         WHEN "010101101010" => data <= X"24FEFF03";
         WHEN "010101101011" => data <= X"004010AA";
         WHEN "010101101100" => data <= X"00F0201A";
         WHEN "010101101101" => data <= X"004031AA";
         WHEN "010101101110" => data <= X"008830E4";
         WHEN "010101101111" => data <= X"08000010";
         WHEN "010101110000" => data <= X"00000015";
         WHEN "010101110001" => data <= X"00F0A018";
         WHEN "010101110010" => data <= X"76FCFF07";
         WHEN "010101110011" => data <= X"421EA59C";
         WHEN "010101110100" => data <= X"0000001B";
         WHEN "010101110101" => data <= X"19FEFF03";
         WHEN "010101110110" => data <= X"0004001A";
         WHEN "010101110111" => data <= X"00F0A018";
         WHEN "010101111000" => data <= X"70FCFF07";
         WHEN "010101111001" => data <= X"551EA59C";
         WHEN "010101111010" => data <= X"0000001B";
         WHEN "010101111011" => data <= X"13FEFF03";
         WHEN "010101111100" => data <= X"0000001A";
         WHEN "010101111101" => data <= X"00007084";
         WHEN "010101111110" => data <= X"D3FDFF07";
         WHEN "010101111111" => data <= X"00000015";
         WHEN "010110000000" => data <= X"0000201A";
         WHEN "010110000001" => data <= X"00880BE4";
         WHEN "010110000010" => data <= X"05000010";
         WHEN "010110000011" => data <= X"3F00201A";
         WHEN "010110000100" => data <= X"00F0A018";
         WHEN "010110000101" => data <= X"ADFEFF03";
         WHEN "010110000110" => data <= X"8A1EA59C";
         WHEN "010110000111" => data <= X"FFFF31AA";
         WHEN "010110001000" => data <= X"04007086";
         WHEN "010110001001" => data <= X"0088B3E4";
         WHEN "010110001010" => data <= X"23000010";
         WHEN "010110001011" => data <= X"0000401B";
         WHEN "010110001100" => data <= X"00F0A018";
         WHEN "010110001101" => data <= X"A5FEFF03";
         WHEN "010110001110" => data <= X"A71EA59C";
         WHEN "010110001111" => data <= X"0088BAE2";
         WHEN "010110010000" => data <= X"00007587";
         WHEN "010110010001" => data <= X"00003A87";
         WHEN "010110010010" => data <= X"00C81BE4";
         WHEN "010110010011" => data <= X"11000010";
         WHEN "010110010100" => data <= X"04883AE2";
         WHEN "010110010101" => data <= X"00F06018";
         WHEN "010110010110" => data <= X"0000B586";
         WHEN "010110010111" => data <= X"04E09CE0";
         WHEN "010110011000" => data <= X"00003A87";
         WHEN "010110011001" => data <= X"180B639C";
         WHEN "010110011010" => data <= X"08C801D4";
         WHEN "010110011011" => data <= X"04A801D4";
         WHEN "010110011100" => data <= X"008801D4";
         WHEN "010110011101" => data <= X"18B801D4";
         WHEN "010110011110" => data <= X"149801D4";
         WHEN "010110011111" => data <= X"49FCFF07";
         WHEN "010110100000" => data <= X"0C2801D4";
         WHEN "010110100001" => data <= X"1800E186";
         WHEN "010110100010" => data <= X"14006186";
         WHEN "010110100011" => data <= X"0C00A184";
         WHEN "010110100100" => data <= X"0100739E";
         WHEN "010110100101" => data <= X"04005A9F";
         WHEN "010110100110" => data <= X"00003786";
         WHEN "010110100111" => data <= X"009851E4";
         WHEN "010110101000" => data <= X"E7FFFF13";
         WHEN "010110101001" => data <= X"0004201A";
         WHEN "010110101010" => data <= X"00F0A018";
         WHEN "010110101011" => data <= X"87FEFF03";
         WHEN "010110101100" => data <= X"ED1EA59C";
         WHEN "010110101101" => data <= X"00F0A018";
         WHEN "010110101110" => data <= X"00F0801B";
         WHEN "010110101111" => data <= X"0000601A";
         WHEN "010110110000" => data <= X"0400E0AA";
         WHEN "010110110001" => data <= X"C71EA59C";
         WHEN "010110110010" => data <= X"F4FFFF03";
         WHEN "010110110011" => data <= X"B0099C9F";
         WHEN "010110110100" => data <= X"00F0201A";
         WHEN "010110110101" => data <= X"004031AA";
         WHEN "010110110110" => data <= X"00F0801B";
         WHEN "010110110111" => data <= X"00F0401B";
         WHEN "010110111000" => data <= X"008810E4";
         WHEN "010110111001" => data <= X"B0099C9F";
         WHEN "010110111010" => data <= X"06000010";
         WHEN "010110111011" => data <= X"180B5A9F";
         WHEN "010110111100" => data <= X"0004201A";
         WHEN "010110111101" => data <= X"008830E4";
         WHEN "010110111110" => data <= X"07000010";
         WHEN "010110111111" => data <= X"00000015";
         WHEN "010111000000" => data <= X"00F0A018";
         WHEN "010111000001" => data <= X"681EA59C";
         WHEN "010111000010" => data <= X"04E09CE0";
         WHEN "010111000011" => data <= X"73FEFF03";
         WHEN "010111000100" => data <= X"04D07AE0";
         WHEN "010111000101" => data <= X"00007084";
         WHEN "010111000110" => data <= X"8BFDFF07";
         WHEN "010111000111" => data <= X"00000015";
         WHEN "010111001000" => data <= X"0000201A";
         WHEN "010111001001" => data <= X"00880BE4";
         WHEN "010111001010" => data <= X"05000010";
         WHEN "010111001011" => data <= X"3F00201A";
         WHEN "010111001100" => data <= X"00F0A018";
         WHEN "010111001101" => data <= X"F5FFFF03";
         WHEN "010111001110" => data <= X"8A1EA59C";
         WHEN "010111001111" => data <= X"FFFF31AA";
         WHEN "010111010000" => data <= X"04007086";
         WHEN "010111010001" => data <= X"0088B3E4";
         WHEN "010111010010" => data <= X"04000010";
         WHEN "010111010011" => data <= X"00F0A018";
         WHEN "010111010100" => data <= X"EEFFFF03";
         WHEN "010111010101" => data <= X"A71EA59C";
         WHEN "010111010110" => data <= X"00F0A018";
         WHEN "010111010111" => data <= X"FB1EA59C";
         WHEN "010111011000" => data <= X"04E09CE0";
         WHEN "010111011001" => data <= X"0FFCFF07";
         WHEN "010111011010" => data <= X"04D07AE0";
         WHEN "010111011011" => data <= X"00F0A018";
         WHEN "010111011100" => data <= X"0004201A";
         WHEN "010111011101" => data <= X"0000601A";
         WHEN "010111011110" => data <= X"FFFFE0AE";
         WHEN "010111011111" => data <= X"00FC201B";
         WHEN "010111100000" => data <= X"1E1FA59C";
         WHEN "010111100001" => data <= X"0400A0AA";
         WHEN "010111100010" => data <= X"0000B586";
         WHEN "010111100011" => data <= X"009855E4";
         WHEN "010111100100" => data <= X"0E000010";
         WHEN "010111100101" => data <= X"04E09CE0";
         WHEN "010111100110" => data <= X"00F0A018";
         WHEN "010111100111" => data <= X"451FA59C";
         WHEN "010111101000" => data <= X"00FCFF07";
         WHEN "010111101001" => data <= X"04D07AE0";
         WHEN "010111101010" => data <= X"040020AA";
         WHEN "010111101011" => data <= X"00006018";
         WHEN "010111101100" => data <= X"00009184";
         WHEN "010111101101" => data <= X"FCFAFF07";
         WHEN "010111101110" => data <= X"00000015";
         WHEN "010111101111" => data <= X"00F0A018";
         WHEN "010111110000" => data <= X"D2FFFF03";
         WHEN "010111110001" => data <= X"5E1FA59C";
         WHEN "010111110010" => data <= X"0000B186";
         WHEN "010111110011" => data <= X"00B815E4";
         WHEN "010111110100" => data <= X"14000010";
         WHEN "010111110101" => data <= X"00C8B1E2";
         WHEN "010111110110" => data <= X"00A801D4";
         WHEN "010111110111" => data <= X"04E09CE0";
         WHEN "010111111000" => data <= X"04D07AE0";
         WHEN "010111111001" => data <= X"28B801D4";
         WHEN "010111111010" => data <= X"249801D4";
         WHEN "010111111011" => data <= X"20C801D4";
         WHEN "010111111100" => data <= X"188801D4";
         WHEN "010111111101" => data <= X"0C2801D4";
         WHEN "010111111110" => data <= X"EAFBFF07";
         WHEN "010111111111" => data <= X"14A801D4";
         WHEN "011000000000" => data <= X"1400A186";
         WHEN "011000000001" => data <= X"E1FAFF07";
         WHEN "011000000010" => data <= X"04A875E0";
         WHEN "011000000011" => data <= X"2800E186";
         WHEN "011000000100" => data <= X"24006186";
         WHEN "011000000101" => data <= X"20002187";
         WHEN "011000000110" => data <= X"18002186";
         WHEN "011000000111" => data <= X"0C00A184";
         WHEN "011000001000" => data <= X"0100739E";
         WHEN "011000001001" => data <= X"D8FFFF03";
         WHEN "011000001010" => data <= X"0400319E";
         WHEN "011000001011" => data <= X"00F0801B";
         WHEN "011000001100" => data <= X"00F0401B";
         WHEN "011000001101" => data <= X"B0099C9F";
         WHEN "011000001110" => data <= X"180B5A9F";
         WHEN "011000001111" => data <= X"00F0A018";
         WHEN "011000010000" => data <= X"741FA59C";
         WHEN "011000010001" => data <= X"04E09CE0";
         WHEN "011000010010" => data <= X"D6FBFF07";
         WHEN "011000010011" => data <= X"04D07AE0";
         WHEN "011000010100" => data <= X"00F0A018";
         WHEN "011000010101" => data <= X"0004201A";
         WHEN "011000010110" => data <= X"FFFFE0AE";
         WHEN "011000010111" => data <= X"00FC201B";
         WHEN "011000011000" => data <= X"1E1FA59C";
         WHEN "011000011001" => data <= X"0005A01A";
         WHEN "011000011010" => data <= X"00007186";
         WHEN "011000011011" => data <= X"00B813E4";
         WHEN "011000011100" => data <= X"14000010";
         WHEN "011000011101" => data <= X"00C871E2";
         WHEN "011000011110" => data <= X"009801D4";
         WHEN "011000011111" => data <= X"04E09CE0";
         WHEN "011000100000" => data <= X"04D07AE0";
         WHEN "011000100001" => data <= X"28A801D4";
         WHEN "011000100010" => data <= X"24B801D4";
         WHEN "011000100011" => data <= X"20C801D4";
         WHEN "011000100100" => data <= X"188801D4";
         WHEN "011000100101" => data <= X"0C2801D4";
         WHEN "011000100110" => data <= X"C2FBFF07";
         WHEN "011000100111" => data <= X"149801D4";
         WHEN "011000101000" => data <= X"14006186";
         WHEN "011000101001" => data <= X"B9FAFF07";
         WHEN "011000101010" => data <= X"049873E0";
         WHEN "011000101011" => data <= X"2800A186";
         WHEN "011000101100" => data <= X"2400E186";
         WHEN "011000101101" => data <= X"20002187";
         WHEN "011000101110" => data <= X"18002186";
         WHEN "011000101111" => data <= X"0C00A184";
         WHEN "011000110000" => data <= X"0400319E";
         WHEN "011000110001" => data <= X"00A831E4";
         WHEN "011000110010" => data <= X"E8FFFF13";
         WHEN "011000110011" => data <= X"00000015";
         WHEN "011000110100" => data <= X"00F0A018";
         WHEN "011000110101" => data <= X"8DFFFF03";
         WHEN "011000110110" => data <= X"921FA59C";
         WHEN "011000110111" => data <= X"0100189F";
         WHEN "011000111000" => data <= X"008838E4";
         WHEN "011000111001" => data <= X"66FEFF13";
         WHEN "011000111010" => data <= X"04D09AE0";
         WHEN "011000111011" => data <= X"A5FEFF03";
         WHEN "011000111100" => data <= X"00F0A018";
         WHEN "011000111101" => data <= X"00F0A018";
         WHEN "011000111110" => data <= X"AAFBFF07";
         WHEN "011000111111" => data <= X"4F20A59C";
         WHEN "011001000000" => data <= X"4EFDFF03";
         WHEN "011001000001" => data <= X"04D0DAE3";
         WHEN "011001000010" => data <= X"39FCFF07";
         WHEN "011001000011" => data <= X"270080AB";
         WHEN "011001000100" => data <= X"37FCFF07";
         WHEN "011001000101" => data <= X"FF004BA7";
         WHEN "011001000110" => data <= X"D0FF5A9F";
         WHEN "011001000111" => data <= X"020020AA";
         WHEN "011001001000" => data <= X"08883AE2";
         WHEN "011001001001" => data <= X"FF004BA6";
         WHEN "011001001010" => data <= X"00D031E2";
         WHEN "011001001011" => data <= X"008831E2";
         WHEN "011001001100" => data <= X"D0FF529E";
         WHEN "011001001101" => data <= X"42FDFF03";
         WHEN "011001001110" => data <= X"008852E2";
         WHEN "011001001111" => data <= X"6720A59C";
         WHEN "011001010000" => data <= X"E4FDFF03";
         WHEN "011001010001" => data <= X"00008018";
         WHEN "011001010010" => data <= X"1A000010";
         WHEN "011001010011" => data <= X"080020AA";
         WHEN "011001010100" => data <= X"0888D6E2";
         WHEN "011001010101" => data <= X"0100CE9D";
         WHEN "011001010110" => data <= X"040020AA";
         WHEN "011001010111" => data <= X"00882EE4";
         WHEN "011001011000" => data <= X"48000010";
         WHEN "011001011001" => data <= X"00B0DCE2";
         WHEN "011001011010" => data <= X"10002186";
         WHEN "011001011011" => data <= X"008830E4";
         WHEN "011001011100" => data <= X"17000010";
         WHEN "011001011101" => data <= X"0004201A";
         WHEN "011001011110" => data <= X"FF0F20AA";
         WHEN "011001011111" => data <= X"008834E4";
         WHEN "011001100000" => data <= X"0E000010";
         WHEN "011001100001" => data <= X"008854E4";
         WHEN "011001100010" => data <= X"00F0A018";
         WHEN "011001100011" => data <= X"00F08018";
         WHEN "011001100100" => data <= X"00F06018";
         WHEN "011001100101" => data <= X"7520A59C";
         WHEN "011001100110" => data <= X"B009849C";
         WHEN "011001100111" => data <= X"81FBFF07";
         WHEN "011001101000" => data <= X"180B639C";
         WHEN "011001101001" => data <= X"010040AA";
         WHEN "011001101010" => data <= X"07000000";
         WHEN "011001101011" => data <= X"001080AA";
         WHEN "011001101100" => data <= X"E9FFFF03";
         WHEN "011001101101" => data <= X"0000C01A";
         WHEN "011001101110" => data <= X"1500000C";
         WHEN "011001101111" => data <= X"020020AA";
         WHEN "011001110000" => data <= X"010040AA";
         WHEN "011001110001" => data <= X"1DFDFF03";
         WHEN "011001110010" => data <= X"0000001B";
         WHEN "011001110011" => data <= X"008830E4";
         WHEN "011001110100" => data <= X"0F000010";
         WHEN "011001110101" => data <= X"020020AA";
         WHEN "011001110110" => data <= X"0000201A";
         WHEN "011001110111" => data <= X"008834E4";
         WHEN "011001111000" => data <= X"16FDFF13";
         WHEN "011001111001" => data <= X"010040AA";
         WHEN "011001111010" => data <= X"00F0A018";
         WHEN "011001111011" => data <= X"00F08018";
         WHEN "011001111100" => data <= X"00F06018";
         WHEN "011001111101" => data <= X"A420A59C";
         WHEN "011001111110" => data <= X"B009849C";
         WHEN "011001111111" => data <= X"69FBFF07";
         WHEN "011010000000" => data <= X"180B639C";
         WHEN "011010000001" => data <= X"0DFDFF03";
         WHEN "011010000010" => data <= X"049092E2";
         WHEN "011010000011" => data <= X"0888D4E1";
         WHEN "011010000100" => data <= X"0000601A";
         WHEN "011010000101" => data <= X"FF3F34A6";
         WHEN "011010000110" => data <= X"009831E4";
         WHEN "011010000111" => data <= X"08000010";
         WHEN "011010001000" => data <= X"00F0A018";
         WHEN "011010001001" => data <= X"00F06018";
         WHEN "011010001010" => data <= X"007001D4";
         WHEN "011010001011" => data <= X"C520A59C";
         WHEN "011010001100" => data <= X"00008018";
         WHEN "011010001101" => data <= X"5BFBFF07";
         WHEN "011010001110" => data <= X"180B639C";
         WHEN "011010001111" => data <= X"0000201A";
         WHEN "011010010000" => data <= X"008802E4";
         WHEN "011010010001" => data <= X"11000010";
         WHEN "011010010010" => data <= X"007030E2";
         WHEN "011010010011" => data <= X"01007672";
         WHEN "011010010100" => data <= X"009811D4";
         WHEN "011010010101" => data <= X"0100949E";
         WHEN "011010010110" => data <= X"00A078E4";
         WHEN "011010010111" => data <= X"09000010";
         WHEN "011010011000" => data <= X"0000C019";
         WHEN "011010011001" => data <= X"0000201A";
         WHEN "011010011010" => data <= X"008802E4";
         WHEN "011010011011" => data <= X"03000010";
         WHEN "011010011100" => data <= X"00000015";
         WHEN "011010011101" => data <= X"04A010D4";
         WHEN "011010011110" => data <= X"04A014E3";
         WHEN "011010011111" => data <= X"0000C019";
         WHEN "011010100000" => data <= X"70FDFF03";
         WHEN "011010100001" => data <= X"FFFF529E";
         WHEN "011010100010" => data <= X"00003186";
         WHEN "011010100011" => data <= X"01003172";
         WHEN "011010100100" => data <= X"008816E4";
         WHEN "011010100101" => data <= X"F0FFFF13";
         WHEN "011010100110" => data <= X"04D0BAE0";
         WHEN "011010100111" => data <= X"00F06018";
         WHEN "011010101000" => data <= X"08B001D4";
         WHEN "011010101001" => data <= X"048801D4";
         WHEN "011010101010" => data <= X"007001D4";
         WHEN "011010101011" => data <= X"00008018";
         WHEN "011010101100" => data <= X"3CFBFF07";
         WHEN "011010101101" => data <= X"180B639C";
         WHEN "011010101110" => data <= X"E8FFFF03";
         WHEN "011010101111" => data <= X"0100949E";
         WHEN "011010110000" => data <= X"20737562";
         WHEN "011010110001" => data <= X"6F727265";
         WHEN "011010110010" => data <= X"000A2172";
         WHEN "011010110011" => data <= X"61746144";
         WHEN "011010110100" => data <= X"67617020";
         WHEN "011010110101" => data <= X"61662065";
         WHEN "011010110110" => data <= X"0A746C75";
         WHEN "011010110111" => data <= X"70206900";
         WHEN "011010111000" => data <= X"20656761";
         WHEN "011010111001" => data <= X"6C756166";
         WHEN "011010111010" => data <= X"74000A74";
         WHEN "011010111011" => data <= X"0A6B6369";
         WHEN "011010111100" => data <= X"6C6C6100";
         WHEN "011010111101" => data <= X"216E6769";
         WHEN "011010111110" => data <= X"3F3F000A";
         WHEN "011010111111" => data <= X"000A3F3F";
         WHEN "011011000000" => data <= X"676E6970";
         WHEN "011011000001" => data <= X"7464000A";
         WHEN "011011000010" => data <= X"000A626C";
         WHEN "011011000011" => data <= X"626C7469";
         WHEN "011011000100" => data <= X"6152000A";
         WHEN "011011000101" => data <= X"2165676E";
         WHEN "011011000110" => data <= X"7953000A";
         WHEN "011011000111" => data <= X"6C616373";
         WHEN "011011001000" => data <= X"54000A6C";
         WHEN "011011001001" => data <= X"21706172";
         WHEN "011011001010" => data <= X"7242000A";
         WHEN "011011001011" => data <= X"0A6B6165";
         WHEN "011011001100" => data <= X"65684300";
         WHEN "011011001101" => data <= X"6E696B63";
         WHEN "011011001110" => data <= X"616C2067";
         WHEN "011011001111" => data <= X"70207473";
         WHEN "011011010000" => data <= X"20656761";
         WHEN "011011010001" => data <= X"6620666F";
         WHEN "011011010010" => data <= X"6873616C";
         WHEN "011011010011" => data <= X"706D6520";
         WHEN "011011010100" => data <= X"000A7974";
         WHEN "011011010101" => data <= X"73616C46";
         WHEN "011011010110" => data <= X"72652068";
         WHEN "011011010111" => data <= X"21726F72";
         WHEN "011011011000" => data <= X"7245000A";
         WHEN "011011011001" => data <= X"6E697361";
         WHEN "011011011010" => data <= X"616C2067";
         WHEN "011011011011" => data <= X"70207473";
         WHEN "011011011100" => data <= X"20656761";
         WHEN "011011011101" => data <= X"4620666F";
         WHEN "011011011110" => data <= X"6873616C";
         WHEN "011011011111" => data <= X"7257000A";
         WHEN "011011100000" => data <= X"6E697469";
         WHEN "011011100001" => data <= X"65742067";
         WHEN "011011100010" => data <= X"73207473";
         WHEN "011011100011" => data <= X"65757165";
         WHEN "011011100100" => data <= X"2065636E";
         WHEN "011011100101" => data <= X"66206F74";
         WHEN "011011100110" => data <= X"6873616C";
         WHEN "011011100111" => data <= X"56000A2E";
         WHEN "011011101000" => data <= X"66697265";
         WHEN "011011101001" => data <= X"676E6979";
         WHEN "011011101010" => data <= X"73657420";
         WHEN "011011101011" => data <= X"65732074";
         WHEN "011011101100" => data <= X"6E657571";
         WHEN "011011101101" => data <= X"66206563";
         WHEN "011011101110" => data <= X"206D6F72";
         WHEN "011011101111" => data <= X"73616C66";
         WHEN "011011110000" => data <= X"000A2E68";
         WHEN "011011110001" => data <= X"74736554";
         WHEN "011011110010" => data <= X"69616620";
         WHEN "011011110011" => data <= X"3A64656C";
         WHEN "011011110100" => data <= X"20642520";
         WHEN "011011110101" => data <= X"7830203A";
         WHEN "011011110110" => data <= X"2F205825";
         WHEN "011011110111" => data <= X"7830203D";
         WHEN "011011111000" => data <= X"000A5825";
         WHEN "011011111001" => data <= X"73616C46";
         WHEN "011011111010" => data <= X"65742068";
         WHEN "011011111011" => data <= X"6F207473";
         WHEN "011011111100" => data <= X"2E79616B";
         WHEN "011011111101" => data <= X"43000A0A";
         WHEN "011011111110" => data <= X"37342D53";
         WHEN "011011111111" => data <= X"79532033";
         WHEN "011100000000" => data <= X"6D657473";
         WHEN "011100000001" => data <= X"6F727020";
         WHEN "011100000010" => data <= X"6D617267";
         WHEN "011100000011" => data <= X"676E696D";
         WHEN "011100000100" => data <= X"726F6620";
         WHEN "011100000101" => data <= X"73797320";
         WHEN "011100000110" => data <= X"736D6574";
         WHEN "011100000111" => data <= X"206E6F20";
         WHEN "011100001000" => data <= X"70696863";
         WHEN "011100001001" => data <= X"704F000A";
         WHEN "011100001010" => data <= X"69726E65";
         WHEN "011100001011" => data <= X"62206373";
         WHEN "011100001100" => data <= X"64657361";
         WHEN "011100001101" => data <= X"72697620";
         WHEN "011100001110" => data <= X"6C617574";
         WHEN "011100001111" => data <= X"6F725020";
         WHEN "011100010000" => data <= X"79746F74";
         WHEN "011100010001" => data <= X"0A2E6570";
         WHEN "011100010010" => data <= X"69754200";
         WHEN "011100010011" => data <= X"7620646C";
         WHEN "011100010100" => data <= X"69737265";
         WHEN "011100010101" => data <= X"203A6E6F";
         WHEN "011100010110" => data <= X"206E6F4D";
         WHEN "011100010111" => data <= X"20706553";
         WHEN "011100011000" => data <= X"31203220";
         WHEN "011100011001" => data <= X"39353A30";
         WHEN "011100011010" => data <= X"2032303A";
         WHEN "011100011011" => data <= X"43204D41";
         WHEN "011100011100" => data <= X"20545345";
         WHEN "011100011101" => data <= X"34323032";
         WHEN "011100011110" => data <= X"49000A0A";
         WHEN "011100011111" => data <= X"206D6120";
         WHEN "011100100000" => data <= X"20555043";
         WHEN "011100100001" => data <= X"6F206425";
         WHEN "011100100010" => data <= X"64252066";
         WHEN "011100100011" => data <= X"6E757220";
         WHEN "011100100100" => data <= X"676E696E";
         WHEN "011100100101" => data <= X"20746120";
         WHEN "011100100110" => data <= X"25642500";
         WHEN "011100100111" => data <= X"64252E64";
         WHEN "011100101000" => data <= X"4D206425";
         WHEN "011100101001" => data <= X"0A2E7A48";
         WHEN "011100101010" => data <= X"6157000A";
         WHEN "011100101011" => data <= X"6E697469";
         WHEN "011100101100" => data <= X"6F662067";
         WHEN "011100101101" => data <= X"50432072";
         WHEN "011100101110" => data <= X"20312055";
         WHEN "011100101111" => data <= X"61206F74";
         WHEN "011100110000" => data <= X"76697463";
         WHEN "011100110001" => data <= X"20657461";
         WHEN "011100110010" => data <= X"000A656D";
         WHEN "011100110011" => data <= X"706D754A";
         WHEN "011100110100" => data <= X"20676E69";
         WHEN "011100110101" => data <= X"6D206F74";
         WHEN "011100110110" => data <= X"206E6961";
         WHEN "011100110111" => data <= X"676F7270";
         WHEN "011100111000" => data <= X"206D6172";
         WHEN "011100111001" => data <= X"25783040";
         WHEN "011100111010" => data <= X"50000A58";
         WHEN "011100111011" => data <= X"72676F72";
         WHEN "011100111100" => data <= X"70206D61";
         WHEN "011100111101" => data <= X"65736572";
         WHEN "011100111110" => data <= X"6220746E";
         WHEN "011100111111" => data <= X"6E207475";
         WHEN "011101000000" => data <= X"6620746F";
         WHEN "011101000001" => data <= X"7420726F";
         WHEN "011101000010" => data <= X"20736968";
         WHEN "011101000011" => data <= X"67726154";
         WHEN "011101000100" => data <= X"0A2E7465";
         WHEN "011101000101" => data <= X"20646944";
         WHEN "011101000110" => data <= X"20756F79";
         WHEN "011101000111" => data <= X"6F6C7075";
         WHEN "011101001000" => data <= X"66206461";
         WHEN "011101001001" => data <= X"7420726F";
         WHEN "011101001010" => data <= X"4F206568";
         WHEN "011101001011" => data <= X"32343152";
         WHEN "011101001100" => data <= X"6C702030";
         WHEN "011101001101" => data <= X"6F667461";
         WHEN "011101001110" => data <= X"0A3F6D72";
         WHEN "011101001111" => data <= X"776F4400";
         WHEN "011101010000" => data <= X"616F6C6E";
         WHEN "011101010001" => data <= X"64203A64";
         WHEN "011101010010" => data <= X"0A656E6F";
         WHEN "011101010011" => data <= X"61655200";
         WHEN "011101010100" => data <= X"676E6964";
         WHEN "011101010101" => data <= X"646F6320";
         WHEN "011101010110" => data <= X"61742065";
         WHEN "011101010111" => data <= X"0A656C62";
         WHEN "011101011000" => data <= X"776F4400";
         WHEN "011101011001" => data <= X"616F6C6E";
         WHEN "011101011010" => data <= X"73203A64";
         WHEN "011101011011" => data <= X"61207465";
         WHEN "011101011100" => data <= X"65726464";
         WHEN "011101011101" => data <= X"3D207373";
         WHEN "011101011110" => data <= X"25783020";
         WHEN "011101011111" => data <= X"45000A58";
         WHEN "011101100000" => data <= X"726F7272";
         WHEN "011101100001" => data <= X"6F6E202C";
         WHEN "011101100010" => data <= X"6F727020";
         WHEN "011101100011" => data <= X"6D617267";
         WHEN "011101100100" => data <= X"616F6C20";
         WHEN "011101100101" => data <= X"21646564";
         WHEN "011101100110" => data <= X"754A000A";
         WHEN "011101100111" => data <= X"6E69706D";
         WHEN "011101101000" => data <= X"6F742067";
         WHEN "011101101001" => data <= X"6F727020";
         WHEN "011101101010" => data <= X"6D617267";
         WHEN "011101101011" => data <= X"45000A6D";
         WHEN "011101101100" => data <= X"726F7272";
         WHEN "011101101101" => data <= X"6F6E202C";
         WHEN "011101101110" => data <= X"6F727020";
         WHEN "011101101111" => data <= X"6D617267";
         WHEN "011101110000" => data <= X"206E6920";
         WHEN "011101110001" => data <= X"73616C46";
         WHEN "011101110010" => data <= X"000A2168";
         WHEN "011101110011" => data <= X"74746553";
         WHEN "011101110100" => data <= X"20676E69";
         WHEN "011101110101" => data <= X"676F7270";
         WHEN "011101110110" => data <= X"6F6D202E";
         WHEN "011101110111" => data <= X"000A6564";
         WHEN "011101111000" => data <= X"74746553";
         WHEN "011101111001" => data <= X"20676E69";
         WHEN "011101111010" => data <= X"69726576";
         WHEN "011101111011" => data <= X"6D202E66";
         WHEN "011101111100" => data <= X"0A65646F";
         WHEN "011101111101" => data <= X"206F4E00";
         WHEN "011101111110" => data <= X"676F7270";
         WHEN "011101111111" => data <= X"206D6172";
         WHEN "011110000000" => data <= X"73657270";
         WHEN "011110000001" => data <= X"0A746E65";
         WHEN "011110000010" => data <= X"6F725000";
         WHEN "011110000011" => data <= X"6D617267";
         WHEN "011110000100" => data <= X"206E6920";
         WHEN "011110000101" => data <= X"206D656D";
         WHEN "011110000110" => data <= X"6D6F7266";
         WHEN "011110000111" => data <= X"25783020";
         WHEN "011110001000" => data <= X"6F742058";
         WHEN "011110001001" => data <= X"25783020";
         WHEN "011110001010" => data <= X"53000A58";
         WHEN "011110001011" => data <= X"63746977";
         WHEN "011110001100" => data <= X"20646568";
         WHEN "011110001101" => data <= X"73206F74";
         WHEN "011110001110" => data <= X"2D74666F";
         WHEN "011110001111" => data <= X"736F6962";
         WHEN "011110010000" => data <= X"7753000A";
         WHEN "011110010001" => data <= X"68637469";
         WHEN "011110010010" => data <= X"74206465";
         WHEN "011110010011" => data <= X"6C46206F";
         WHEN "011110010100" => data <= X"0A687361";
         WHEN "011110010101" => data <= X"69775300";
         WHEN "011110010110" => data <= X"65686374";
         WHEN "011110010111" => data <= X"6F742064";
         WHEN "011110011000" => data <= X"52445320";
         WHEN "011110011001" => data <= X"000A6D61";
         WHEN "011110011010" => data <= X"61656C50";
         WHEN "011110011011" => data <= X"63206573";
         WHEN "011110011100" => data <= X"676E6168";
         WHEN "011110011101" => data <= X"6F742065";
         WHEN "011110011110" => data <= X"65687420";
         WHEN "011110011111" => data <= X"52445320";
         WHEN "011110100000" => data <= X"62204D41";
         WHEN "011110100001" => data <= X"742A2079";
         WHEN "011110100010" => data <= X"6F4E000A";
         WHEN "011110100011" => data <= X"6F727020";
         WHEN "011110100100" => data <= X"6D617267";
         WHEN "011110100101" => data <= X"616F6C20";
         WHEN "011110100110" => data <= X"20646564";
         WHEN "011110100111" => data <= X"53206E69";
         WHEN "011110101000" => data <= X"6D615244";
         WHEN "011110101001" => data <= X"50000A21";
         WHEN "011110101010" => data <= X"72676F72";
         WHEN "011110101011" => data <= X"64206D61";
         WHEN "011110101100" => data <= X"2073656F";
         WHEN "011110101101" => data <= X"20746F6E";
         WHEN "011110101110" => data <= X"20746966";
         WHEN "011110101111" => data <= X"46206E69";
         WHEN "011110110000" => data <= X"6873616C";
         WHEN "011110110001" => data <= X"43000A21";
         WHEN "011110110010" => data <= X"61706D6F";
         WHEN "011110110011" => data <= X"65206572";
         WHEN "011110110100" => data <= X"726F7272";
         WHEN "011110110101" => data <= X"20746120";
         WHEN "011110110110" => data <= X"58257830";
         WHEN "011110110111" => data <= X"30203A20";
         WHEN "011110111000" => data <= X"20582578";
         WHEN "011110111001" => data <= X"30203D21";
         WHEN "011110111010" => data <= X"0A582578";
         WHEN "011110111011" => data <= X"6D6F4300";
         WHEN "011110111100" => data <= X"65726170";
         WHEN "011110111101" => data <= X"6E6F6420";
         WHEN "011110111110" => data <= X"43000A65";
         WHEN "011110111111" => data <= X"6B636568";
         WHEN "011111000000" => data <= X"20676E69";
         WHEN "011111000001" => data <= X"74206669";
         WHEN "011111000010" => data <= X"66206568";
         WHEN "011111000011" => data <= X"6873616C";
         WHEN "011111000100" => data <= X"20736920";
         WHEN "011111000101" => data <= X"74706D65";
         WHEN "011111000110" => data <= X"2E2E2E79";
         WHEN "011111000111" => data <= X"7453000A";
         WHEN "011111001000" => data <= X"20747261";
         WHEN "011111001001" => data <= X"73616C66";
         WHEN "011111001010" => data <= X"72652068";
         WHEN "011111001011" => data <= X"20657361";
         WHEN "011111001100" => data <= X"6C637963";
         WHEN "011111001101" => data <= X"6F662065";
         WHEN "011111001110" => data <= X"61702072";
         WHEN "011111001111" => data <= X"30206567";
         WHEN "011111010000" => data <= X"0A582578";
         WHEN "011111010001" => data <= X"61745300";
         WHEN "011111010010" => data <= X"70207472";
         WHEN "011111010011" => data <= X"72676F72";
         WHEN "011111010100" => data <= X"696D6D61";
         WHEN "011111010101" => data <= X"6620676E";
         WHEN "011111010110" => data <= X"6873616C";
         WHEN "011111010111" => data <= X"7250000A";
         WHEN "011111011000" => data <= X"6172676F";
         WHEN "011111011001" => data <= X"6E696D6D";
         WHEN "011111011010" => data <= X"69662067";
         WHEN "011111011011" => data <= X"6873696E";
         WHEN "011111011100" => data <= X"000A6465";
         WHEN "011111011101" => data <= X"63656843";
         WHEN "011111011110" => data <= X"676E696B";
         WHEN "011111011111" => data <= X"20666920";
         WHEN "011111100000" => data <= X"73616C66";
         WHEN "011111100001" => data <= X"73692068";
         WHEN "011111100010" => data <= X"69642720";
         WHEN "011111100011" => data <= X"27797472";
         WHEN "011111100100" => data <= X"6C46000A";
         WHEN "011111100101" => data <= X"20687361";
         WHEN "011111100110" => data <= X"65207369";
         WHEN "011111100111" => data <= X"7974706D";
         WHEN "011111101000" => data <= X"72652820";
         WHEN "011111101001" => data <= X"64657361";
         WHEN "011111101010" => data <= X"0A0A2E29";
         WHEN "011111101011" => data <= X"61745300";
         WHEN "011111101100" => data <= X"6E697472";
         WHEN "011111101101" => data <= X"69732067";
         WHEN "011111101110" => data <= X"656C706D";
         WHEN "011111101111" => data <= X"52445320";
         WHEN "011111110000" => data <= X"6D206D61";
         WHEN "011111110001" => data <= X"68636D65";
         WHEN "011111110010" => data <= X"2E6B6365";
         WHEN "011111110011" => data <= X"57000A0A";
         WHEN "011111110100" => data <= X"69746972";
         WHEN "011111110101" => data <= X"2E2E676E";
         WHEN "011111110110" => data <= X"56000A2E";
         WHEN "011111110111" => data <= X"66697265";
         WHEN "011111111000" => data <= X"676E6979";
         WHEN "011111111001" => data <= X"0A2E2E2E";
         WHEN "011111111010" => data <= X"72724500";
         WHEN "011111111011" => data <= X"4020726F";
         WHEN "011111111100" => data <= X"58257830";
         WHEN "011111111101" => data <= X"30203A20";
         WHEN "011111111110" => data <= X"20582578";
         WHEN "011111111111" => data <= X"30203D21";
         WHEN "100000000000" => data <= X"0A582578";
         WHEN "100000000001" => data <= X"20724E00";
         WHEN "100000000010" => data <= X"6520666F";
         WHEN "100000000011" => data <= X"726F7272";
         WHEN "100000000100" => data <= X"6F662073";
         WHEN "100000000101" => data <= X"20646E75";
         WHEN "100000000110" => data <= X"6425203A";
         WHEN "100000000111" => data <= X"654D000A";
         WHEN "100000001000" => data <= X"6568636D";
         WHEN "100000001001" => data <= X"64206B63";
         WHEN "100000001010" => data <= X"2C656E6F";
         WHEN "100000001011" => data <= X"20642520";
         WHEN "100000001100" => data <= X"6F727265";
         WHEN "100000001101" => data <= X"0A0A7372";
         WHEN "100000001110" => data <= X"74655300";
         WHEN "100000001111" => data <= X"676E6974";
         WHEN "100000010000" => data <= X"61747320";
         WHEN "100000010001" => data <= X"74206B63";
         WHEN "100000010010" => data <= X"5053206F";
         WHEN "100000010011" => data <= X"53000A4D";
         WHEN "100000010100" => data <= X"69747465";
         WHEN "100000010101" => data <= X"7320676E";
         WHEN "100000010110" => data <= X"6B636174";
         WHEN "100000010111" => data <= X"206F7420";
         WHEN "100000011000" => data <= X"41524453";
         WHEN "100000011001" => data <= X"55000A4D";
         WHEN "100000011010" => data <= X"6F6E6B6E";
         WHEN "100000011011" => data <= X"63206E77";
         WHEN "100000011100" => data <= X"2165646F";
         WHEN "100000011101" => data <= X"6F725000";
         WHEN "100000011110" => data <= X"6D617267";
         WHEN "100000011111" => data <= X"6F6F7420";
         WHEN "100000100000" => data <= X"67696220";
         WHEN "100000100001" => data <= X"206F7420";
         WHEN "100000100010" => data <= X"20746966";
         WHEN "100000100011" => data <= X"53206E69";
         WHEN "100000100100" => data <= X"6274666F";
         WHEN "100000100101" => data <= X"2C736F69";
         WHEN "100000100110" => data <= X"6F626120";
         WHEN "100000100111" => data <= X"6E697472";
         WHEN "100000101000" => data <= X"000A2167";
         WHEN "100000101001" => data <= X"6E6E6143";
         WHEN "100000101010" => data <= X"7020746F";
         WHEN "100000101011" => data <= X"72676F72";
         WHEN "100000101100" => data <= X"66206D61";
         WHEN "100000101101" => data <= X"6873616C";
         WHEN "100000101110" => data <= X"6261202C";
         WHEN "100000101111" => data <= X"6974726F";
         WHEN "100000110000" => data <= X"0A21676E";
         WHEN "100000110001" => data <= X"776F4400";
         WHEN "100000110010" => data <= X"616F6C6E";
         WHEN "100000110011" => data <= X"61203A64";
         WHEN "100000110100" => data <= X"78302074";
         WHEN "100000110101" => data <= X"000A5825";
         WHEN "100000110110" => data <= X"69726556";
         WHEN "100000110111" => data <= X"61636966";
         WHEN "100000111000" => data <= X"6E6F6974";
         WHEN "100000111001" => data <= X"72726520";
         WHEN "100000111010" => data <= X"6120726F";
         WHEN "100000111011" => data <= X"78302074";
         WHEN "100000111100" => data <= X"3A205825";
         WHEN "100000111101" => data <= X"25783020";
         WHEN "100000111110" => data <= X"3D212058";
         WHEN "100000111111" => data <= X"25783020";
         WHEN "100001000000" => data <= X"4B000A58";
         WHEN "100001000001" => data <= X"6E776F6E";
         WHEN "100001000010" => data <= X"32535220";
         WHEN "100001000011" => data <= X"63203233";
         WHEN "100001000100" => data <= X"616D6D6F";
         WHEN "100001000101" => data <= X"3A73646E";
         WHEN "100001000110" => data <= X"2024000A";
         WHEN "100001000111" => data <= X"61745320";
         WHEN "100001001000" => data <= X"74207472";
         WHEN "100001001001" => data <= X"70206568";
         WHEN "100001001010" => data <= X"72676F72";
         WHEN "100001001011" => data <= X"6C206D61";
         WHEN "100001001100" => data <= X"6564616F";
         WHEN "100001001101" => data <= X"6E692064";
         WHEN "100001001110" => data <= X"72617420";
         WHEN "100001001111" => data <= X"0A746567";
         WHEN "100001010000" => data <= X"20702A00";
         WHEN "100001010001" => data <= X"20746553";
         WHEN "100001010010" => data <= X"676F7270";
         WHEN "100001010011" => data <= X"6D6D6172";
         WHEN "100001010100" => data <= X"20676E69";
         WHEN "100001010101" => data <= X"65646F6D";
         WHEN "100001010110" => data <= X"65642820";
         WHEN "100001010111" => data <= X"6C756166";
         WHEN "100001011000" => data <= X"000A2974";
         WHEN "100001011001" => data <= X"5320762A";
         WHEN "100001011010" => data <= X"76207465";
         WHEN "100001011011" => data <= X"66697265";
         WHEN "100001011100" => data <= X"74616369";
         WHEN "100001011101" => data <= X"206E6F69";
         WHEN "100001011110" => data <= X"65646F6D";
         WHEN "100001011111" => data <= X"692A000A";
         WHEN "100001100000" => data <= X"6F685320";
         WHEN "100001100001" => data <= X"6E692077";
         WHEN "100001100010" => data <= X"6F206F66";
         WHEN "100001100011" => data <= X"7270206E";
         WHEN "100001100100" => data <= X"6172676F";
         WHEN "100001100101" => data <= X"6E69206D";
         WHEN "100001100110" => data <= X"72617420";
         WHEN "100001100111" => data <= X"0A746567";
         WHEN "100001101000" => data <= X"20742A00";
         WHEN "100001101001" => data <= X"67676F54";
         WHEN "100001101010" => data <= X"7420656C";
         WHEN "100001101011" => data <= X"65677261";
         WHEN "100001101100" => data <= X"65622074";
         WHEN "100001101101" => data <= X"65657774";
         WHEN "100001101110" => data <= X"4453206E";
         WHEN "100001101111" => data <= X"206D6152";
         WHEN "100001110000" => data <= X"66656428";
         WHEN "100001110001" => data <= X"746C7561";
         WHEN "100001110010" => data <= X"73202C29";
         WHEN "100001110011" => data <= X"2D74666F";
         WHEN "100001110100" => data <= X"736F6942";
         WHEN "100001110101" => data <= X"646E6120";
         WHEN "100001110110" => data <= X"616C4620";
         WHEN "100001110111" => data <= X"000A6873";
         WHEN "100001111000" => data <= X"50206D2A";
         WHEN "100001111001" => data <= X"6F667265";
         WHEN "100001111010" => data <= X"73206D72";
         WHEN "100001111011" => data <= X"6C706D69";
         WHEN "100001111100" => data <= X"44532065";
         WHEN "100001111101" => data <= X"206D6152";
         WHEN "100001111110" => data <= X"636D656D";
         WHEN "100001111111" => data <= X"6B636568";
         WHEN "100010000000" => data <= X"732A000A";
         WHEN "100010000001" => data <= X"65684320";
         WHEN "100010000010" => data <= X"53206B63";
         WHEN "100010000011" => data <= X"662D4950";
         WHEN "100010000100" => data <= X"6873616C";
         WHEN "100010000101" => data <= X"69686320";
         WHEN "100010000110" => data <= X"2A000A70";
         WHEN "100010000111" => data <= X"72452065";
         WHEN "100010001000" => data <= X"20657361";
         WHEN "100010001001" => data <= X"2D495053";
         WHEN "100010001010" => data <= X"73616C46";
         WHEN "100010001011" => data <= X"68632068";
         WHEN "100010001100" => data <= X"000A7069";
         WHEN "100010001101" => data <= X"5320662A";
         WHEN "100010001110" => data <= X"65726F74";
         WHEN "100010001111" => data <= X"6F727020";
         WHEN "100010010000" => data <= X"6D617267";
         WHEN "100010010001" => data <= X"616F6C20";
         WHEN "100010010010" => data <= X"20646564";
         WHEN "100010010011" => data <= X"53206E69";
         WHEN "100010010100" => data <= X"4D415244";
         WHEN "100010010101" => data <= X"206F7420";
         WHEN "100010010110" => data <= X"2D495053";
         WHEN "100010010111" => data <= X"73616C46";
         WHEN "100010011000" => data <= X"2A000A68";
         WHEN "100010011001" => data <= X"6F432063";
         WHEN "100010011010" => data <= X"7261706D";
         WHEN "100010011011" => data <= X"72702065";
         WHEN "100010011100" => data <= X"6172676F";
         WHEN "100010011101" => data <= X"6F6C206D";
         WHEN "100010011110" => data <= X"64656461";
         WHEN "100010011111" => data <= X"206E6920";
         WHEN "100010100000" => data <= X"41524453";
         WHEN "100010100001" => data <= X"6977204D";
         WHEN "100010100010" => data <= X"53206874";
         WHEN "100010100011" => data <= X"462D4950";
         WHEN "100010100100" => data <= X"6873616C";
         WHEN "100010100101" => data <= X"722A000A";
         WHEN "100010100110" => data <= X"6E755220";
         WHEN "100010100111" => data <= X"6F727020";
         WHEN "100010101000" => data <= X"6D617267";
         WHEN "100010101001" => data <= X"6F747320";
         WHEN "100010101010" => data <= X"20646572";
         WHEN "100010101011" => data <= X"53206E69";
         WHEN "100010101100" => data <= X"462D4950";
         WHEN "100010101101" => data <= X"6873616C";
         WHEN "100010101110" => data <= X"712A000A";
         WHEN "100010101111" => data <= X"676F5420";
         WHEN "100010110000" => data <= X"20656C67";
         WHEN "100010110001" => data <= X"63617473";
         WHEN "100010110010" => data <= X"6F70206B";
         WHEN "100010110011" => data <= X"65746E69";
         WHEN "100010110100" => data <= X"72662072";
         WHEN "100010110101" => data <= X"53206D6F";
         WHEN "100010110110" => data <= X"4D415244";
         WHEN "100010110111" => data <= X"65642820";
         WHEN "100010111000" => data <= X"6C756166";
         WHEN "100010111001" => data <= X"77202974";
         WHEN "100010111010" => data <= X"20687469";
         WHEN "100010111011" => data <= X"0A4D5053";
         WHEN "100010111100" => data <= X"20682A00";
         WHEN "100010111101" => data <= X"73696854";
         WHEN "100010111110" => data <= X"6C656820";
         WHEN "100010111111" => data <= X"72637370";
         WHEN "100011000000" => data <= X"0A6E6565";
         WHEN "100011000001" => data <= X"0000000A";
         WHEN "100011000010" => data <= X"EFBEADDE";
         WHEN "100011000011" => data <= X"01000000";
         WHEN "100011000100" => data <= X"02000000";
         WHEN "100011000101" => data <= X"03000000";
         WHEN "100011000110" => data <= X"04000000";
         WHEN "100011000111" => data <= X"05000000";
         WHEN "100011001000" => data <= X"06000000";
         WHEN "100011001001" => data <= X"07000000";
         WHEN "100011001010" => data <= X"032100F0";
         WHEN "100011001011" => data <= X"1A2100F0";
         WHEN "100011001100" => data <= X"412100F0";
         WHEN "100011001101" => data <= X"642100F0";
         WHEN "100011001110" => data <= X"7E2100F0";
         WHEN "100011001111" => data <= X"A12100F0";
         WHEN "100011010000" => data <= X"E02100F0";
         WHEN "100011010001" => data <= X"022200F0";
         WHEN "100011010010" => data <= X"1B2200F0";
         WHEN "100011010011" => data <= X"342200F0";
         WHEN "100011010100" => data <= X"632200F0";
         WHEN "100011010101" => data <= X"962200F0";
         WHEN "100011010110" => data <= X"BA2200F0";
         WHEN "100011010111" => data <= X"F12200F0";
         WHEN OTHERS => data <= X"00000000";
      END CASE;
   END PROCESS TheRom;

END platform_independent;

--------------------------------------------------------------------------------
-- $RCSfile: $
--
-- DESC    : OpenRisk 1420 
--
-- AUTHOR  : Dr. Theo Kluter
--
-- CVS     : $Revision: $
--           $Date: $
--           $Author: $
--           $Source: $
--
--------------------------------------------------------------------------------
--
--  HISTORY :
--
--  $Log: 
--------------------------------------------------------------------------------

ARCHITECTURE platform_independent OF bios_rom IS

BEGIN

   TheRom : PROCESS( address )
   BEGIN
      CASE (address) IS
         WHEN "00000000000" => data <= X"2014ADDE";
         WHEN "00000000001" => data <= X"00000015";
         WHEN "00000000010" => data <= X"11000000";
         WHEN "00000000011" => data <= X"00000015";
         WHEN "00000000100" => data <= X"0F000000";
         WHEN "00000000101" => data <= X"00000015";
         WHEN "00000000110" => data <= X"0D000000";
         WHEN "00000000111" => data <= X"00000015";
         WHEN "00000001000" => data <= X"0B000000";
         WHEN "00000001001" => data <= X"00000015";
         WHEN "00000001010" => data <= X"09000000";
         WHEN "00000001011" => data <= X"00000015";
         WHEN "00000001100" => data <= X"00C02018";
         WHEN "00000001101" => data <= X"FC1F21A8";
         WHEN "00000001110" => data <= X"050060E0";
         WHEN "00000001111" => data <= X"0C030004";
         WHEN "00000010000" => data <= X"050080E0";
         WHEN "00000010010" => data <= X"00000015";
         WHEN "00000010011" => data <= X"84FF219C";
         WHEN "00000010100" => data <= X"001001D4";
         WHEN "00000010101" => data <= X"041801D4";
         WHEN "00000010110" => data <= X"082001D4";
         WHEN "00000010111" => data <= X"0C2801D4";
         WHEN "00000011000" => data <= X"103001D4";
         WHEN "00000011001" => data <= X"143801D4";
         WHEN "00000011010" => data <= X"184001D4";
         WHEN "00000011011" => data <= X"1C4801D4";
         WHEN "00000011100" => data <= X"205001D4";
         WHEN "00000011101" => data <= X"245801D4";
         WHEN "00000011110" => data <= X"286001D4";
         WHEN "00000011111" => data <= X"2C6801D4";
         WHEN "00000100000" => data <= X"307001D4";
         WHEN "00000100001" => data <= X"347801D4";
         WHEN "00000100010" => data <= X"388001D4";
         WHEN "00000100011" => data <= X"3C8801D4";
         WHEN "00000100100" => data <= X"409001D4";
         WHEN "00000100101" => data <= X"449801D4";
         WHEN "00000100110" => data <= X"48A001D4";
         WHEN "00000100111" => data <= X"4CA801D4";
         WHEN "00000101000" => data <= X"50B001D4";
         WHEN "00000101001" => data <= X"54B801D4";
         WHEN "00000101010" => data <= X"58C001D4";
         WHEN "00000101011" => data <= X"5CC801D4";
         WHEN "00000101100" => data <= X"60D001D4";
         WHEN "00000101101" => data <= X"64D801D4";
         WHEN "00000101110" => data <= X"68E001D4";
         WHEN "00000101111" => data <= X"6CE801D4";
         WHEN "00000110000" => data <= X"70F001D4";
         WHEN "00000110001" => data <= X"74F801D4";
         WHEN "00000110010" => data <= X"1200E0B7";
         WHEN "00000110011" => data <= X"0200FFBB";
         WHEN "00000110100" => data <= X"00F0C01B";
         WHEN "00000110101" => data <= X"6C01DEAB";
         WHEN "00000110110" => data <= X"00F8DEE3";
         WHEN "00000110111" => data <= X"0000FE87";
         WHEN "00000111000" => data <= X"00F80048";
         WHEN "00000111001" => data <= X"00000015";
         WHEN "00000111010" => data <= X"00004184";
         WHEN "00000111011" => data <= X"04006184";
         WHEN "00000111100" => data <= X"08008184";
         WHEN "00000111101" => data <= X"0C00A184";
         WHEN "00000111110" => data <= X"1000C184";
         WHEN "00000111111" => data <= X"1400E184";
         WHEN "00001000000" => data <= X"18000185";
         WHEN "00001000001" => data <= X"1C002185";
         WHEN "00001000010" => data <= X"20004185";
         WHEN "00001000011" => data <= X"24006185";
         WHEN "00001000100" => data <= X"28008185";
         WHEN "00001000101" => data <= X"2C00A185";
         WHEN "00001000110" => data <= X"3000C185";
         WHEN "00001000111" => data <= X"3400E185";
         WHEN "00001001000" => data <= X"38000186";
         WHEN "00001001001" => data <= X"3C002186";
         WHEN "00001001010" => data <= X"40004186";
         WHEN "00001001011" => data <= X"44006186";
         WHEN "00001001100" => data <= X"48008186";
         WHEN "00001001101" => data <= X"4C00A186";
         WHEN "00001001110" => data <= X"5000C186";
         WHEN "00001001111" => data <= X"5400E186";
         WHEN "00001010000" => data <= X"58000187";
         WHEN "00001010001" => data <= X"5C002187";
         WHEN "00001010010" => data <= X"60004187";
         WHEN "00001010011" => data <= X"64006187";
         WHEN "00001010100" => data <= X"68008187";
         WHEN "00001010101" => data <= X"6C00A187";
         WHEN "00001010110" => data <= X"7000C187";
         WHEN "00001010111" => data <= X"7400E187";
         WHEN "00001011000" => data <= X"7C00219C";
         WHEN "00001011001" => data <= X"00000024";
         WHEN "00001011010" => data <= X"00000015";
         WHEN "00001011011" => data <= X"300000F0";
         WHEN "00001011100" => data <= X"840100F0";
         WHEN "00001011101" => data <= X"A00100F0";
         WHEN "00001011110" => data <= X"BC0100F0";
         WHEN "00001011111" => data <= X"D80100F0";
         WHEN "00001100000" => data <= X"F40100F0";
         WHEN "00001100001" => data <= X"00F0A018";
         WHEN "00001100010" => data <= X"00F08018";
         WHEN "00001100011" => data <= X"00F06018";
         WHEN "00001100100" => data <= X"6018A59C";
         WHEN "00001100101" => data <= X"8C08849C";
         WHEN "00001100110" => data <= X"39010000";
         WHEN "00001100111" => data <= X"F409639C";
         WHEN "00001101000" => data <= X"00F0A018";
         WHEN "00001101001" => data <= X"00F08018";
         WHEN "00001101010" => data <= X"00F06018";
         WHEN "00001101011" => data <= X"6B18A59C";
         WHEN "00001101100" => data <= X"8C08849C";
         WHEN "00001101101" => data <= X"32010000";
         WHEN "00001101110" => data <= X"F409639C";
         WHEN "00001101111" => data <= X"00F0A018";
         WHEN "00001110000" => data <= X"00F08018";
         WHEN "00001110001" => data <= X"00F06018";
         WHEN "00001110010" => data <= X"7518A59C";
         WHEN "00001110011" => data <= X"8C08849C";
         WHEN "00001110100" => data <= X"2B010000";
         WHEN "00001110101" => data <= X"F409639C";
         WHEN "00001110110" => data <= X"00F0A018";
         WHEN "00001110111" => data <= X"00F08018";
         WHEN "00001111000" => data <= X"00F06018";
         WHEN "00001111001" => data <= X"7A18A59C";
         WHEN "00001111010" => data <= X"8C08849C";
         WHEN "00001111011" => data <= X"24010000";
         WHEN "00001111100" => data <= X"F409639C";
         WHEN "00001111101" => data <= X"00F0A018";
         WHEN "00001111110" => data <= X"00F08018";
         WHEN "00001111111" => data <= X"00F06018";
         WHEN "00010000000" => data <= X"7F18A59C";
         WHEN "00010000001" => data <= X"8C08849C";
         WHEN "00010000010" => data <= X"1D010000";
         WHEN "00010000011" => data <= X"F409639C";
         WHEN "00010000100" => data <= X"0000601A";
         WHEN "00010000101" => data <= X"0700A0AA";
         WHEN "00010000110" => data <= X"02A83372";
         WHEN "00010000111" => data <= X"0000E01A";
         WHEN "00010001000" => data <= X"010031A6";
         WHEN "00010001001" => data <= X"00B831E4";
         WHEN "00010001010" => data <= X"FCFFFF13";
         WHEN "00010001011" => data <= X"00000015";
         WHEN "00010001100" => data <= X"00480044";
         WHEN "00010001101" => data <= X"00000015";
         WHEN "00010001110" => data <= X"00006019";
         WHEN "00010001111" => data <= X"02186B71";
         WHEN "00010010000" => data <= X"00480044";
         WHEN "00010010001" => data <= X"00000015";
         WHEN "00010010010" => data <= X"160020AA";
         WHEN "00010010011" => data <= X"02890370";
         WHEN "00010010100" => data <= X"020020AA";
         WHEN "00010010101" => data <= X"070060AA";
         WHEN "00010010110" => data <= X"02991170";
         WHEN "00010010111" => data <= X"EDFFFF03";
         WHEN "00010011000" => data <= X"00000015";
         WHEN "00010011001" => data <= X"DCFF219C";
         WHEN "00010011010" => data <= X"008001D4";
         WHEN "00010011011" => data <= X"049001D4";
         WHEN "00010011100" => data <= X"08A001D4";
         WHEN "00010011101" => data <= X"0CB001D4";
         WHEN "00010011110" => data <= X"10C001D4";
         WHEN "00010011111" => data <= X"14D001D4";
         WHEN "00010100000" => data <= X"18E001D4";
         WHEN "00010100001" => data <= X"1CF001D4";
         WHEN "00010100010" => data <= X"204801D4";
         WHEN "00010100011" => data <= X"0418C3E2";
         WHEN "00010100100" => data <= X"042044E2";
         WHEN "00010100101" => data <= X"0000001A";
         WHEN "00010100110" => data <= X"0000801A";
         WHEN "00010100111" => data <= X"160000AB";
         WHEN "00010101000" => data <= X"200040AB";
         WHEN "00010101001" => data <= X"010080AB";
         WHEN "00010101010" => data <= X"0700C0AB";
         WHEN "00010101011" => data <= X"009094E5";
         WHEN "00010101100" => data <= X"0C000010";
         WHEN "00010101101" => data <= X"20002185";
         WHEN "00010101110" => data <= X"00000186";
         WHEN "00010101111" => data <= X"04004186";
         WHEN "00010110000" => data <= X"08008186";
         WHEN "00010110001" => data <= X"0C00C186";
         WHEN "00010110010" => data <= X"10000187";
         WHEN "00010110011" => data <= X"14004187";
         WHEN "00010110100" => data <= X"18008187";
         WHEN "00010110101" => data <= X"1C00C187";
         WHEN "00010110110" => data <= X"00480044";
         WHEN "00010110111" => data <= X"2400219C";
         WHEN "00010111000" => data <= X"02C11070";
         WHEN "00010111001" => data <= X"180020AA";
         WHEN "00010111010" => data <= X"008076E2";
         WHEN "00010111011" => data <= X"0000B386";
         WHEN "00010111100" => data <= X"0102B572";
         WHEN "00010111101" => data <= X"02891570";
         WHEN "00010111110" => data <= X"0100319E";
         WHEN "00010111111" => data <= X"00D031E4";
         WHEN "00011000000" => data <= X"FBFFFF13";
         WHEN "00011000001" => data <= X"0400739E";
         WHEN "00011000010" => data <= X"02F11C70";
         WHEN "00011000011" => data <= X"C1FFFF07";
         WHEN "00011000100" => data <= X"0800949E";
         WHEN "00011000101" => data <= X"E6FFFF03";
         WHEN "00011000110" => data <= X"2000109E";
         WHEN "00011000111" => data <= X"B4FF219C";
         WHEN "00011001000" => data <= X"00F08018";
         WHEN "00011001001" => data <= X"2000A0A8";
         WHEN "00011001010" => data <= X"741F849C";
         WHEN "00011001011" => data <= X"0C00619C";
         WHEN "00011001100" => data <= X"2C8001D4";
         WHEN "00011001101" => data <= X"309001D4";
         WHEN "00011001110" => data <= X"38B001D4";
         WHEN "00011001111" => data <= X"3CC001D4";
         WHEN "00011010000" => data <= X"40D001D4";
         WHEN "00011010001" => data <= X"44E001D4";
         WHEN "00011010010" => data <= X"484801D4";
         WHEN "00011010011" => data <= X"34A001D4";
         WHEN "00011010100" => data <= X"AE010004";
         WHEN "00011010101" => data <= X"00F0401A";
         WHEN "00011010110" => data <= X"00F0001A";
         WHEN "00011010111" => data <= X"8C08529E";
         WHEN "00011011000" => data <= X"F409109E";
         WHEN "00011011001" => data <= X"00F0A018";
         WHEN "00011011010" => data <= X"8818A59C";
         WHEN "00011011011" => data <= X"049092E0";
         WHEN "00011011100" => data <= X"C3000004";
         WHEN "00011011101" => data <= X"048070E0";
         WHEN "00011011110" => data <= X"1F00201A";
         WHEN "00011011111" => data <= X"00F0C01A";
         WHEN "00011100000" => data <= X"0000601A";
         WHEN "00011100001" => data <= X"00FC31AA";
         WHEN "00011100010" => data <= X"0004001B";
         WHEN "00011100011" => data <= X"FFFF40AF";
         WHEN "00011100100" => data <= X"B918D69E";
         WHEN "00011100101" => data <= X"010080AB";
         WHEN "00011100110" => data <= X"0200A0AA";
         WHEN "00011100111" => data <= X"08A891E2";
         WHEN "00011101000" => data <= X"00C094E2";
         WHEN "00011101001" => data <= X"0000B486";
         WHEN "00011101010" => data <= X"00D015E4";
         WHEN "00011101011" => data <= X"1D000010";
         WHEN "00011101100" => data <= X"0100319E";
         WHEN "00011101101" => data <= X"0000201A";
         WHEN "00011101110" => data <= X"008813E4";
         WHEN "00011101111" => data <= X"10000010";
         WHEN "00011110000" => data <= X"04B0B6E0";
         WHEN "00011110001" => data <= X"00F0A018";
         WHEN "00011110010" => data <= X"AB18A59C";
         WHEN "00011110011" => data <= X"049092E0";
         WHEN "00011110100" => data <= X"048070E0";
         WHEN "00011110101" => data <= X"30004186";
         WHEN "00011110110" => data <= X"2C000186";
         WHEN "00011110111" => data <= X"34008186";
         WHEN "00011111000" => data <= X"3800C186";
         WHEN "00011111001" => data <= X"3C000187";
         WHEN "00011111010" => data <= X"40004187";
         WHEN "00011111011" => data <= X"44008187";
         WHEN "00011111100" => data <= X"48002185";
         WHEN "00011111101" => data <= X"A2000000";
         WHEN "00011111110" => data <= X"4C00219C";
         WHEN "00011111111" => data <= X"049092E0";
         WHEN "00100000000" => data <= X"9F000004";
         WHEN "00100000001" => data <= X"048070E0";
         WHEN "00100000010" => data <= X"90FFFF07";
         WHEN "00100000011" => data <= X"04A074E0";
         WHEN "00100000100" => data <= X"1F00201A";
         WHEN "00100000101" => data <= X"04E07CE2";
         WHEN "00100000110" => data <= X"00FC31AA";
         WHEN "00100000111" => data <= X"0100319E";
         WHEN "00100001000" => data <= X"2000A01A";
         WHEN "00100001001" => data <= X"00A831E4";
         WHEN "00100001010" => data <= X"DDFFFF13";
         WHEN "00100001011" => data <= X"0200A0AA";
         WHEN "00100001100" => data <= X"00F0A018";
         WHEN "00100001101" => data <= X"D518A59C";
         WHEN "00100001110" => data <= X"049092E0";
         WHEN "00100001111" => data <= X"90000004";
         WHEN "00100010000" => data <= X"048070E0";
         WHEN "00100010001" => data <= X"0C00819E";
         WHEN "00100010010" => data <= X"04A074E2";
         WHEN "00100010011" => data <= X"180020AA";
         WHEN "00100010100" => data <= X"2000E0AA";
         WHEN "00100010101" => data <= X"0000B386";
         WHEN "00100010110" => data <= X"0102B572";
         WHEN "00100010111" => data <= X"02891570";
         WHEN "00100011000" => data <= X"0100319E";
         WHEN "00100011001" => data <= X"00B831E4";
         WHEN "00100011010" => data <= X"FBFFFF13";
         WHEN "00100011011" => data <= X"0400739E";
         WHEN "00100011100" => data <= X"7F00201A";
         WHEN "00100011101" => data <= X"00F031AA";
         WHEN "00100011110" => data <= X"160060AA";
         WHEN "00100011111" => data <= X"02991170";
         WHEN "00100100000" => data <= X"010020AA";
         WHEN "00100100001" => data <= X"070060AA";
         WHEN "00100100010" => data <= X"02991170";
         WHEN "00100100011" => data <= X"61FFFF07";
         WHEN "00100100100" => data <= X"00000015";
         WHEN "00100100101" => data <= X"00F0A018";
         WHEN "00100100110" => data <= X"F618A59C";
         WHEN "00100100111" => data <= X"049092E0";
         WHEN "00100101000" => data <= X"77000004";
         WHEN "00100101001" => data <= X"048070E0";
         WHEN "00100101010" => data <= X"7F04201A";
         WHEN "00100101011" => data <= X"00F031AA";
         WHEN "00100101100" => data <= X"0000601A";
         WHEN "00100101101" => data <= X"080020AB";
         WHEN "00100101110" => data <= X"0000B186";
         WHEN "00100101111" => data <= X"0000F486";
         WHEN "00100110000" => data <= X"00A817E4";
         WHEN "00100110001" => data <= X"14000010";
         WHEN "00100110010" => data <= X"0400319E";
         WHEN "00100110011" => data <= X"00F0A018";
         WHEN "00100110100" => data <= X"08B801D4";
         WHEN "00100110101" => data <= X"04A801D4";
         WHEN "00100110110" => data <= X"009801D4";
         WHEN "00100110111" => data <= X"049092E0";
         WHEN "00100111000" => data <= X"048070E0";
         WHEN "00100111001" => data <= X"66000004";
         WHEN "00100111010" => data <= X"1B19A59C";
         WHEN "00100111011" => data <= X"48002185";
         WHEN "00100111100" => data <= X"2C000186";
         WHEN "00100111101" => data <= X"30004186";
         WHEN "00100111110" => data <= X"34008186";
         WHEN "00100111111" => data <= X"3800C186";
         WHEN "00101000000" => data <= X"3C000187";
         WHEN "00101000001" => data <= X"40004187";
         WHEN "00101000010" => data <= X"44008187";
         WHEN "00101000011" => data <= X"00480044";
         WHEN "00101000100" => data <= X"4C00219C";
         WHEN "00101000101" => data <= X"0100739E";
         WHEN "00101000110" => data <= X"00C833E4";
         WHEN "00101000111" => data <= X"E7FFFF13";
         WHEN "00101001000" => data <= X"0400949E";
         WHEN "00101001001" => data <= X"00F0A018";
         WHEN "00101001010" => data <= X"A9FFFF03";
         WHEN "00101001011" => data <= X"3B19A59C";
         WHEN "00101001100" => data <= X"E8FF219C";
         WHEN "00101001101" => data <= X"008001D4";
         WHEN "00101001110" => data <= X"049001D4";
         WHEN "00101001111" => data <= X"08A001D4";
         WHEN "00101010000" => data <= X"0CB001D4";
         WHEN "00101010001" => data <= X"10C001D4";
         WHEN "00101010010" => data <= X"144801D4";
         WHEN "00101010011" => data <= X"041843E2";
         WHEN "00101010100" => data <= X"042084E2";
         WHEN "00101010101" => data <= X"1C0000AA";
         WHEN "00101010110" => data <= X"090000AB";
         WHEN "00101010111" => data <= X"FCFFC0AE";
         WHEN "00101011000" => data <= X"488074E0";
         WHEN "00101011001" => data <= X"0F0023A6";
         WHEN "00101011010" => data <= X"00C051E4";
         WHEN "00101011011" => data <= X"03000010";
         WHEN "00101011100" => data <= X"3700719C";
         WHEN "00101011101" => data <= X"3000719C";
         WHEN "00101011110" => data <= X"00900048";
         WHEN "00101011111" => data <= X"FCFF109E";
         WHEN "00101100000" => data <= X"00B030E4";
         WHEN "00101100001" => data <= X"F8FFFF13";
         WHEN "00101100010" => data <= X"488074E0";
         WHEN "00101100011" => data <= X"00000186";
         WHEN "00101100100" => data <= X"04004186";
         WHEN "00101100101" => data <= X"08008186";
         WHEN "00101100110" => data <= X"0C00C186";
         WHEN "00101100111" => data <= X"10000187";
         WHEN "00101101000" => data <= X"14002185";
         WHEN "00101101001" => data <= X"00480044";
         WHEN "00101101010" => data <= X"1800219C";
         WHEN "00101101011" => data <= X"DCFF219C";
         WHEN "00101101100" => data <= X"0C8001D4";
         WHEN "00101101101" => data <= X"109001D4";
         WHEN "00101101110" => data <= X"14A001D4";
         WHEN "00101101111" => data <= X"18B001D4";
         WHEN "00101110000" => data <= X"1CC001D4";
         WHEN "00101110001" => data <= X"204801D4";
         WHEN "00101110010" => data <= X"0418C3E2";
         WHEN "00101110011" => data <= X"042044E2";
         WHEN "00101110100" => data <= X"0000801A";
         WHEN "00101110101" => data <= X"0000001A";
         WHEN "00101110110" => data <= X"0A0000AB";
         WHEN "00101110111" => data <= X"04C098E0";
         WHEN "00101111000" => data <= X"9B040004";
         WHEN "00101111001" => data <= X"049072E0";
         WHEN "00101111010" => data <= X"0200219E";
         WHEN "00101111011" => data <= X"00A031E2";
         WHEN "00101111100" => data <= X"30006B9D";
         WHEN "00101111101" => data <= X"005811D8";
         WHEN "00101111110" => data <= X"0000201A";
         WHEN "00101111111" => data <= X"008814E4";
         WHEN "00110000000" => data <= X"04000010";
         WHEN "00110000001" => data <= X"008812E4";
         WHEN "00110000010" => data <= X"05000010";
         WHEN "00110000011" => data <= X"049072E0";
         WHEN "00110000100" => data <= X"0100109E";
         WHEN "00110000101" => data <= X"FF0010A6";
         WHEN "00110000110" => data <= X"049072E0";
         WHEN "00110000111" => data <= X"73040004";
         WHEN "00110001000" => data <= X"04C098E0";
         WHEN "00110001001" => data <= X"0100949E";
         WHEN "00110001010" => data <= X"00C034E4";
         WHEN "00110001011" => data <= X"ECFFFF13";
         WHEN "00110001100" => data <= X"04584BE2";
         WHEN "00110001101" => data <= X"0000201A";
         WHEN "00110001110" => data <= X"008830E4";
         WHEN "00110001111" => data <= X"0A000010";
         WHEN "00110010000" => data <= X"FFFF109E";
         WHEN "00110010001" => data <= X"0C000186";
         WHEN "00110010010" => data <= X"10004186";
         WHEN "00110010011" => data <= X"14008186";
         WHEN "00110010100" => data <= X"1800C186";
         WHEN "00110010101" => data <= X"1C000187";
         WHEN "00110010110" => data <= X"20002185";
         WHEN "00110010111" => data <= X"00480044";
         WHEN "00110011000" => data <= X"2400219C";
         WHEN "00110011001" => data <= X"0200219E";
         WHEN "00110011010" => data <= X"008031E2";
         WHEN "00110011011" => data <= X"00B00048";
         WHEN "00110011100" => data <= X"0000718C";
         WHEN "00110011101" => data <= X"F1FFFF03";
         WHEN "00110011110" => data <= X"0000201A";
         WHEN "00110011111" => data <= X"E0FF219C";
         WHEN "00110100000" => data <= X"008001D4";
         WHEN "00110100001" => data <= X"049001D4";
         WHEN "00110100010" => data <= X"08A001D4";
         WHEN "00110100011" => data <= X"0CB001D4";
         WHEN "00110100100" => data <= X"14D001D4";
         WHEN "00110100101" => data <= X"18E001D4";
         WHEN "00110100110" => data <= X"10C001D4";
         WHEN "00110100111" => data <= X"1C4801D4";
         WHEN "00110101000" => data <= X"041883E2";
         WHEN "00110101001" => data <= X"042004E2";
         WHEN "00110101010" => data <= X"042845E2";
         WHEN "00110101011" => data <= X"2000C19E";
         WHEN "00110101100" => data <= X"250040AB";
         WHEN "00110101101" => data <= X"630080AB";
         WHEN "00110101110" => data <= X"00007290";
         WHEN "00110101111" => data <= X"0000201A";
         WHEN "00110110000" => data <= X"008823E4";
         WHEN "00110110001" => data <= X"3B00000C";
         WHEN "00110110010" => data <= X"00D023E4";
         WHEN "00110110011" => data <= X"5A000010";
         WHEN "00110110100" => data <= X"FF0003A7";
         WHEN "00110110101" => data <= X"01003292";
         WHEN "00110110110" => data <= X"00E011E4";
         WHEN "00110110111" => data <= X"4D000010";
         WHEN "00110111000" => data <= X"00E051E5";
         WHEN "00110111001" => data <= X"1B000010";
         WHEN "00110111010" => data <= X"0000601A";
         WHEN "00110111011" => data <= X"009811E4";
         WHEN "00110111100" => data <= X"28000010";
         WHEN "00110111101" => data <= X"580060AA";
         WHEN "00110111110" => data <= X"009811E4";
         WHEN "00110111111" => data <= X"37000010";
         WHEN "00111000000" => data <= X"0400169F";
         WHEN "00111000001" => data <= X"00A00048";
         WHEN "00111000010" => data <= X"250060A8";
         WHEN "00111000011" => data <= X"0000201A";
         WHEN "00111000100" => data <= X"008810E4";
         WHEN "00111000101" => data <= X"04000010";
         WHEN "00111000110" => data <= X"00000015";
         WHEN "00111000111" => data <= X"00800048";
         WHEN "00111001000" => data <= X"250060A8";
         WHEN "00111001001" => data <= X"0100128F";
         WHEN "00111001010" => data <= X"00A00048";
         WHEN "00111001011" => data <= X"04C078E0";
         WHEN "00111001100" => data <= X"0000201A";
         WHEN "00111001101" => data <= X"008810E4";
         WHEN "00111001110" => data <= X"33000010";
         WHEN "00111001111" => data <= X"00000015";
         WHEN "00111010000" => data <= X"00800048";
         WHEN "00111010001" => data <= X"04C078E0";
         WHEN "00111010010" => data <= X"30000000";
         WHEN "00111010011" => data <= X"0100529E";
         WHEN "00111010100" => data <= X"640060AA";
         WHEN "00111010101" => data <= X"009811E4";
         WHEN "00111010110" => data <= X"EBFFFF0F";
         WHEN "00111010111" => data <= X"0400169F";
         WHEN "00111011000" => data <= X"04A074E0";
         WHEN "00111011001" => data <= X"0000D686";
         WHEN "00111011010" => data <= X"91FFFF07";
         WHEN "00111011011" => data <= X"04B096E0";
         WHEN "00111011100" => data <= X"0000201A";
         WHEN "00111011101" => data <= X"008810E4";
         WHEN "00111011110" => data <= X"22000010";
         WHEN "00111011111" => data <= X"04B096E0";
         WHEN "00111100000" => data <= X"8BFFFF07";
         WHEN "00111100001" => data <= X"048070E0";
         WHEN "00111100010" => data <= X"1F000000";
         WHEN "00111100011" => data <= X"04C0D8E2";
         WHEN "00111100100" => data <= X"00A00048";
         WHEN "00111100101" => data <= X"04D07AE0";
         WHEN "00111100110" => data <= X"0000201A";
         WHEN "00111100111" => data <= X"008810E4";
         WHEN "00111101000" => data <= X"04000010";
         WHEN "00111101001" => data <= X"04D07AE0";
         WHEN "00111101010" => data <= X"00800048";
         WHEN "00111101011" => data <= X"00000015";
         WHEN "00111101100" => data <= X"00000186";
         WHEN "00111101101" => data <= X"04004186";
         WHEN "00111101110" => data <= X"08008186";
         WHEN "00111101111" => data <= X"0C00C186";
         WHEN "00111110000" => data <= X"10000187";
         WHEN "00111110001" => data <= X"14004187";
         WHEN "00111110010" => data <= X"18008187";
         WHEN "00111110011" => data <= X"1C002185";
         WHEN "00111110100" => data <= X"00480044";
         WHEN "00111110101" => data <= X"2000219C";
         WHEN "00111110110" => data <= X"04A074E0";
         WHEN "00111110111" => data <= X"0000D686";
         WHEN "00111111000" => data <= X"54FFFF07";
         WHEN "00111111001" => data <= X"04B096E0";
         WHEN "00111111010" => data <= X"0000201A";
         WHEN "00111111011" => data <= X"008810E4";
         WHEN "00111111100" => data <= X"04000010";
         WHEN "00111111101" => data <= X"04B096E0";
         WHEN "00111111110" => data <= X"4EFFFF07";
         WHEN "00111111111" => data <= X"048070E0";
         WHEN "01000000000" => data <= X"04C0D8E2";
         WHEN "01000000001" => data <= X"0100529E";
         WHEN "01000000010" => data <= X"ACFFFF03";
         WHEN "01000000011" => data <= X"0100529E";
         WHEN "01000000100" => data <= X"0300568E";
         WHEN "01000000101" => data <= X"00A00048";
         WHEN "01000000110" => data <= X"049072E0";
         WHEN "01000000111" => data <= X"0000201A";
         WHEN "01000001000" => data <= X"008810E4";
         WHEN "01000001001" => data <= X"E3FFFF13";
         WHEN "01000001010" => data <= X"049072E0";
         WHEN "01000001011" => data <= X"DFFFFF03";
         WHEN "01000001100" => data <= X"00000015";
         WHEN "01000001101" => data <= X"00A00048";
         WHEN "01000001110" => data <= X"04C078E0";
         WHEN "01000001111" => data <= X"0000201A";
         WHEN "01000010000" => data <= X"008810E4";
         WHEN "01000010001" => data <= X"F1FFFF13";
         WHEN "01000010010" => data <= X"00000015";
         WHEN "01000010011" => data <= X"00800048";
         WHEN "01000010100" => data <= X"04C078E0";
         WHEN "01000010101" => data <= X"99FFFF03";
         WHEN "01000010110" => data <= X"0100529E";
         WHEN "01000010111" => data <= X"0050201A";
         WHEN "01000011000" => data <= X"030071AA";
         WHEN "01000011001" => data <= X"83FFA0AE";
         WHEN "01000011010" => data <= X"00A813D8";
         WHEN "01000011011" => data <= X"1B00A0AA";
         WHEN "01000011100" => data <= X"00A811D8";
         WHEN "01000011101" => data <= X"010031AA";
         WHEN "01000011110" => data <= X"000011D8";
         WHEN "01000011111" => data <= X"030020AA";
         WHEN "01000100000" => data <= X"008813D8";
         WHEN "01000100001" => data <= X"00480044";
         WHEN "01000100010" => data <= X"00000015";
         WHEN "01000100011" => data <= X"0050601A";
         WHEN "01000100100" => data <= X"FF0063A4";
         WHEN "01000100101" => data <= X"0500B3AA";
         WHEN "01000100110" => data <= X"0000358E";
         WHEN "01000100111" => data <= X"400031A6";
         WHEN "01000101000" => data <= X"0000E01A";
         WHEN "01000101001" => data <= X"00B811E4";
         WHEN "01000101010" => data <= X"05000010";
         WHEN "01000101011" => data <= X"00000015";
         WHEN "01000101100" => data <= X"001813D8";
         WHEN "01000101101" => data <= X"00480044";
         WHEN "01000101110" => data <= X"00000015";
         WHEN "01000101111" => data <= X"00000015";
         WHEN "01000110000" => data <= X"F6FFFF03";
         WHEN "01000110001" => data <= X"00000015";
         WHEN "01000110010" => data <= X"0050601A";
         WHEN "01000110011" => data <= X"0500B3AA";
         WHEN "01000110100" => data <= X"0000358E";
         WHEN "01000110101" => data <= X"010031A6";
         WHEN "01000110110" => data <= X"0000E01A";
         WHEN "01000110111" => data <= X"00B811E4";
         WHEN "01000111000" => data <= X"FCFFFF13";
         WHEN "01000111001" => data <= X"00000015";
         WHEN "01000111010" => data <= X"0000738D";
         WHEN "01000111011" => data <= X"00480044";
         WHEN "01000111100" => data <= X"00000015";
         WHEN "01000111101" => data <= X"F0FF219C";
         WHEN "01000111110" => data <= X"FF0063A4";
         WHEN "01000111111" => data <= X"008001D4";
         WHEN "01001000000" => data <= X"D0FF039E";
         WHEN "01001000001" => data <= X"FF0030A6";
         WHEN "01001000010" => data <= X"090060AA";
         WHEN "01001000011" => data <= X"049001D4";
         WHEN "01001000100" => data <= X"08A001D4";
         WHEN "01001000101" => data <= X"009851E4";
         WHEN "01001000110" => data <= X"0800000C";
         WHEN "01001000111" => data <= X"0C4801D4";
         WHEN "01001001000" => data <= X"BFFF239E";
         WHEN "01001001001" => data <= X"FF0031A6";
         WHEN "01001001010" => data <= X"050060AA";
         WHEN "01001001011" => data <= X"009851E4";
         WHEN "01001001100" => data <= X"18000010";
         WHEN "01001001101" => data <= X"C9FF039E";
         WHEN "01001001110" => data <= X"090040AA";
         WHEN "01001001111" => data <= X"050080AA";
         WHEN "01001010000" => data <= X"E2FFFF07";
         WHEN "01001010001" => data <= X"00000015";
         WHEN "01001010010" => data <= X"FF006BA5";
         WHEN "01001010011" => data <= X"D0FF2B9E";
         WHEN "01001010100" => data <= X"FF0071A6";
         WHEN "01001010101" => data <= X"009053E4";
         WHEN "01001010110" => data <= X"04000010";
         WHEN "01001010111" => data <= X"0400A0AA";
         WHEN "01001011000" => data <= X"08A810E2";
         WHEN "01001011001" => data <= X"008011E2";
         WHEN "01001011010" => data <= X"BFFF2B9E";
         WHEN "01001011011" => data <= X"FF0031A6";
         WHEN "01001011100" => data <= X"00A051E4";
         WHEN "01001011101" => data <= X"10000010";
         WHEN "01001011110" => data <= X"9FFF2B9E";
         WHEN "01001011111" => data <= X"040020AA";
         WHEN "01001100000" => data <= X"088810E2";
         WHEN "01001100001" => data <= X"C9FF6B9D";
         WHEN "01001100010" => data <= X"EEFFFF03";
         WHEN "01001100011" => data <= X"00800BE2";
         WHEN "01001100100" => data <= X"9FFF239E";
         WHEN "01001100101" => data <= X"FF0031A6";
         WHEN "01001100110" => data <= X"009851E4";
         WHEN "01001100111" => data <= X"04000010";
         WHEN "01001101000" => data <= X"00000015";
         WHEN "01001101001" => data <= X"E5FFFF03";
         WHEN "01001101010" => data <= X"A9FF039E";
         WHEN "01001101011" => data <= X"E3FFFF03";
         WHEN "01001101100" => data <= X"0000001A";
         WHEN "01001101101" => data <= X"FF0031A6";
         WHEN "01001101110" => data <= X"00A051E4";
         WHEN "01001101111" => data <= X"05000010";
         WHEN "01001110000" => data <= X"040020AA";
         WHEN "01001110001" => data <= X"088810E2";
         WHEN "01001110010" => data <= X"F0FFFF03";
         WHEN "01001110011" => data <= X"A9FF6B9D";
         WHEN "01001110100" => data <= X"0090B3E4";
         WHEN "01001110101" => data <= X"DBFFFF13";
         WHEN "01001110110" => data <= X"048070E1";
         WHEN "01001110111" => data <= X"04004186";
         WHEN "01001111000" => data <= X"00000186";
         WHEN "01001111001" => data <= X"08008186";
         WHEN "01001111010" => data <= X"0C002185";
         WHEN "01001111011" => data <= X"00480044";
         WHEN "01001111100" => data <= X"1000219C";
         WHEN "01001111101" => data <= X"FF0063A4";
         WHEN "01001111110" => data <= X"020020AA";
         WHEN "01001111111" => data <= X"00191170";
         WHEN "01010000000" => data <= X"00480044";
         WHEN "01010000001" => data <= X"00000015";
         WHEN "01010000010" => data <= X"041863E1";
         WHEN "01010000011" => data <= X"0000201A";
         WHEN "01010000100" => data <= X"002831E4";
         WHEN "01010000101" => data <= X"04000010";
         WHEN "01010000110" => data <= X"008864E2";
         WHEN "01010000111" => data <= X"00480044";
         WHEN "01010001000" => data <= X"00000015";
         WHEN "01010001001" => data <= X"0000B392";
         WHEN "01010001010" => data <= X"00886BE2";
         WHEN "01010001011" => data <= X"00A813D8";
         WHEN "01010001100" => data <= X"F8FFFF03";
         WHEN "01010001101" => data <= X"0100319E";
         WHEN "01010001110" => data <= X"A8FF219C";
         WHEN "01010001111" => data <= X"00F08018";
         WHEN "01010010000" => data <= X"3800A0A8";
         WHEN "01010010001" => data <= X"941F849C";
         WHEN "01010010010" => data <= X"488001D4";
         WHEN "01010010011" => data <= X"4C9001D4";
         WHEN "01010010100" => data <= X"50A001D4";
         WHEN "01010010101" => data <= X"544801D4";
         WHEN "01010010110" => data <= X"ECFFFF07";
         WHEN "01010010111" => data <= X"1000619C";
         WHEN "01010011000" => data <= X"030020AA";
         WHEN "01010011001" => data <= X"00011170";
         WHEN "01010011010" => data <= X"00F0401A";
         WHEN "01010011011" => data <= X"00F0801A";
         WHEN "01010011100" => data <= X"8C08529E";
         WHEN "01010011101" => data <= X"F409949E";
         WHEN "01010011110" => data <= X"00F0A018";
         WHEN "01010011111" => data <= X"4E19A59C";
         WHEN "01010100000" => data <= X"049092E0";
         WHEN "01010100001" => data <= X"FEFEFF07";
         WHEN "01010100010" => data <= X"04A074E0";
         WHEN "01010100011" => data <= X"00F0A018";
         WHEN "01010100100" => data <= X"6D19A59C";
         WHEN "01010100101" => data <= X"049092E0";
         WHEN "01010100110" => data <= X"F9FEFF07";
         WHEN "01010100111" => data <= X"04A074E0";
         WHEN "01010101000" => data <= X"00F0A018";
         WHEN "01010101001" => data <= X"9019A59C";
         WHEN "01010101010" => data <= X"049092E0";
         WHEN "01010101011" => data <= X"F4FEFF07";
         WHEN "01010101100" => data <= X"04A074E0";
         WHEN "01010101101" => data <= X"FF00201A";
         WHEN "01010101110" => data <= X"FFFF31AA";
         WHEN "01010101111" => data <= X"04000072";
         WHEN "01010110000" => data <= X"0000A01A";
         WHEN "01010110001" => data <= X"038870E2";
         WHEN "01010110010" => data <= X"00A813E4";
         WHEN "01010110011" => data <= X"FCFFFF13";
         WHEN "01010110100" => data <= X"00F0A018";
         WHEN "01010110101" => data <= X"040020AA";
         WHEN "01010110110" => data <= X"488830E2";
         WHEN "01010110111" => data <= X"070031A6";
         WHEN "01010111000" => data <= X"048801D4";
         WHEN "01010111001" => data <= X"070030A6";
         WHEN "01010111010" => data <= X"008801D4";
         WHEN "01010111011" => data <= X"C219A59C";
         WHEN "01010111100" => data <= X"049092E0";
         WHEN "01010111101" => data <= X"E2FEFF07";
         WHEN "01010111110" => data <= X"04A074E0";
         WHEN "01010111111" => data <= X"0C0020AA";
         WHEN "01011000000" => data <= X"488830E2";
         WHEN "01011000001" => data <= X"0F0031A6";
         WHEN "01011000010" => data <= X"0C8801D4";
         WHEN "01011000011" => data <= X"100020AA";
         WHEN "01011000100" => data <= X"488830E2";
         WHEN "01011000101" => data <= X"0F0031A6";
         WHEN "01011000110" => data <= X"088801D4";
         WHEN "01011000111" => data <= X"140020AA";
         WHEN "01011001000" => data <= X"488830E2";
         WHEN "01011001001" => data <= X"0F0031A6";
         WHEN "01011001010" => data <= X"048801D4";
         WHEN "01011001011" => data <= X"180020AA";
         WHEN "01011001100" => data <= X"488830E2";
         WHEN "01011001101" => data <= X"0F0031A6";
         WHEN "01011001110" => data <= X"00F0A018";
         WHEN "01011001111" => data <= X"008801D4";
         WHEN "01011010000" => data <= X"E019A59C";
         WHEN "01011010001" => data <= X"049092E0";
         WHEN "01011010010" => data <= X"CDFEFF07";
         WHEN "01011010011" => data <= X"04A074E0";
         WHEN "01011010100" => data <= X"ADDE201A";
         WHEN "01011010101" => data <= X"0004601A";
         WHEN "01011010110" => data <= X"201431AA";
         WHEN "01011010111" => data <= X"0000B386";
         WHEN "01011011000" => data <= X"008835E4";
         WHEN "01011011001" => data <= X"13000010";
         WHEN "01011011010" => data <= X"0000201A";
         WHEN "01011011011" => data <= X"080010A6";
         WHEN "01011011100" => data <= X"008830E4";
         WHEN "01011011101" => data <= X"0F000010";
         WHEN "01011011110" => data <= X"040033AA";
         WHEN "01011011111" => data <= X"0200A0AA";
         WHEN "01011100000" => data <= X"00003186";
         WHEN "01011100001" => data <= X"08A831E2";
         WHEN "01011100010" => data <= X"008830E4";
         WHEN "01011100011" => data <= X"15000010";
         WHEN "01011100100" => data <= X"0080B3E2";
         WHEN "01011100101" => data <= X"00F0A018";
         WHEN "01011100110" => data <= X"F119A59C";
         WHEN "01011100111" => data <= X"049092E0";
         WHEN "01011101000" => data <= X"B7FEFF07";
         WHEN "01011101001" => data <= X"04A074E0";
         WHEN "01011101010" => data <= X"30000074";
         WHEN "01011101011" => data <= X"00000015";
         WHEN "01011101100" => data <= X"1000019E";
         WHEN "01011101101" => data <= X"0000201A";
         WHEN "01011101110" => data <= X"0000B084";
         WHEN "01011101111" => data <= X"008825E4";
         WHEN "01011110000" => data <= X"0D000010";
         WHEN "01011110001" => data <= X"0400109E";
         WHEN "01011110010" => data <= X"48000186";
         WHEN "01011110011" => data <= X"4C004186";
         WHEN "01011110100" => data <= X"50008186";
         WHEN "01011110101" => data <= X"54002185";
         WHEN "01011110110" => data <= X"00480044";
         WHEN "01011110111" => data <= X"5800219C";
         WHEN "01011111000" => data <= X"0000B586";
         WHEN "01011111001" => data <= X"0400109E";
         WHEN "01011111010" => data <= X"FCAFF0D7";
         WHEN "01011111011" => data <= X"E8FFFF03";
         WHEN "01011111100" => data <= X"008830E4";
         WHEN "01011111101" => data <= X"049092E0";
         WHEN "01011111110" => data <= X"A1FEFF07";
         WHEN "01011111111" => data <= X"04A074E0";
         WHEN "01100000000" => data <= X"EEFFFF03";
         WHEN "01100000001" => data <= X"0000201A";
         WHEN "01100000010" => data <= X"ADDE201A";
         WHEN "01100000011" => data <= X"201471AA";
         WHEN "01100000100" => data <= X"009803E4";
         WHEN "01100000101" => data <= X"13000010";
         WHEN "01100000110" => data <= X"FFFF601A";
         WHEN "01100000111" => data <= X"039863E0";
         WHEN "01100001000" => data <= X"008823E4";
         WHEN "01100001001" => data <= X"10000010";
         WHEN "01100001010" => data <= X"FFFF60AD";
         WHEN "01100001011" => data <= X"00F0A018";
         WHEN "01100001100" => data <= X"00F08018";
         WHEN "01100001101" => data <= X"00F06018";
         WHEN "01100001110" => data <= X"FCFF219C";
         WHEN "01100001111" => data <= X"0D1AA59C";
         WHEN "01100010000" => data <= X"8C08849C";
         WHEN "01100010001" => data <= X"004801D4";
         WHEN "01100010010" => data <= X"8DFEFF07";
         WHEN "01100010011" => data <= X"F409639C";
         WHEN "01100010100" => data <= X"FFFF60AD";
         WHEN "01100010101" => data <= X"00002185";
         WHEN "01100010110" => data <= X"00480044";
         WHEN "01100010111" => data <= X"0400219C";
         WHEN "01100011000" => data <= X"00006019";
         WHEN "01100011001" => data <= X"00480044";
         WHEN "01100011010" => data <= X"00000015";
         WHEN "01100011011" => data <= X"ACFC219C";
         WHEN "01100011100" => data <= X"287301D4";
         WHEN "01100011101" => data <= X"2C8301D4";
         WHEN "01100011110" => data <= X"309301D4";
         WHEN "01100011111" => data <= X"44E301D4";
         WHEN "01100100000" => data <= X"48F301D4";
         WHEN "01100100001" => data <= X"504B01D4";
         WHEN "01100100010" => data <= X"34A301D4";
         WHEN "01100100011" => data <= X"38B301D4";
         WHEN "01100100100" => data <= X"3CC301D4";
         WHEN "01100100101" => data <= X"40D301D4";
         WHEN "01100100110" => data <= X"F1FEFF07";
         WHEN "01100100111" => data <= X"4C1301D4";
         WHEN "01100101000" => data <= X"66FFFF07";
         WHEN "01100101001" => data <= X"010040AA";
         WHEN "01100101010" => data <= X"00F0201A";
         WHEN "01100101011" => data <= X"FC1C319E";
         WHEN "01100101100" => data <= X"0000801B";
         WHEN "01100101101" => data <= X"0000C019";
         WHEN "01100101110" => data <= X"0490D2E3";
         WHEN "01100101111" => data <= X"0000001A";
         WHEN "01100110000" => data <= X"108801D4";
         WHEN "01100110001" => data <= X"270040AB";
         WHEN "01100110010" => data <= X"00FFFF07";
         WHEN "01100110011" => data <= X"00000015";
         WHEN "01100110100" => data <= X"FF000BA7";
         WHEN "01100110101" => data <= X"00D018E4";
         WHEN "01100110110" => data <= X"6F020010";
         WHEN "01100110111" => data <= X"00D058E4";
         WHEN "01100111000" => data <= X"48000010";
         WHEN "01100111001" => data <= X"240020AA";
         WHEN "01100111010" => data <= X"008818E4";
         WHEN "01100111011" => data <= X"9F000010";
         WHEN "01100111100" => data <= X"008858E4";
         WHEN "01100111101" => data <= X"13000010";
         WHEN "01100111110" => data <= X"230020AA";
         WHEN "01100111111" => data <= X"008818E4";
         WHEN "01101000000" => data <= X"93000010";
         WHEN "01101000001" => data <= X"F6FF789E";
         WHEN "01101000010" => data <= X"FF0073A6";
         WHEN "01101000011" => data <= X"160020AA";
         WHEN "01101000100" => data <= X"008853E4";
         WHEN "01101000101" => data <= X"09000010";
         WHEN "01101000110" => data <= X"BFFF201A";
         WHEN "01101000111" => data <= X"F6FF31AA";
         WHEN "01101001000" => data <= X"889831E2";
         WHEN "01101001001" => data <= X"010031A6";
         WHEN "01101001010" => data <= X"0000601A";
         WHEN "01101001011" => data <= X"009831E4";
         WHEN "01101001100" => data <= X"E6FFFF0F";
         WHEN "01101001101" => data <= X"00000015";
         WHEN "01101001110" => data <= X"44000000";
         WHEN "01101001111" => data <= X"00006019";
         WHEN "01101010000" => data <= X"260020AA";
         WHEN "01101010001" => data <= X"008818E4";
         WHEN "01101010010" => data <= X"FCFFFF0F";
         WHEN "01101010011" => data <= X"250000AB";
         WHEN "01101010100" => data <= X"DEFEFF07";
         WHEN "01101010101" => data <= X"0000401B";
         WHEN "01101010110" => data <= X"00F0A018";
         WHEN "01101010111" => data <= X"00F06018";
         WHEN "01101011000" => data <= X"6F1AA59C";
         WHEN "01101011001" => data <= X"00008018";
         WHEN "01101011010" => data <= X"F409639C";
         WHEN "01101011011" => data <= X"44FEFF07";
         WHEN "01101011100" => data <= X"FF004BA4";
         WHEN "01101011101" => data <= X"200000AB";
         WHEN "01101011110" => data <= X"00C002E4";
         WHEN "01101011111" => data <= X"1D000010";
         WHEN "01101100000" => data <= X"00D03AE2";
         WHEN "01101100001" => data <= X"00D031E2";
         WHEN "01101100010" => data <= X"2800619E";
         WHEN "01101100011" => data <= X"0088F3E2";
         WHEN "01101100100" => data <= X"0000A01A";
         WHEN "01101100101" => data <= X"0100B59E";
         WHEN "01101100110" => data <= X"001017D8";
         WHEN "01101100111" => data <= X"188801D4";
         WHEN "01101101000" => data <= X"14A801D4";
         WHEN "01101101001" => data <= X"C9FEFF07";
         WHEN "01101101010" => data <= X"0CB801D4";
         WHEN "01101101011" => data <= X"FF004BA4";
         WHEN "01101101100" => data <= X"00C022E4";
         WHEN "01101101101" => data <= X"0C00E186";
         WHEN "01101101110" => data <= X"1400A186";
         WHEN "01101101111" => data <= X"0100F79E";
         WHEN "01101110000" => data <= X"F5FFFF13";
         WHEN "01101110001" => data <= X"18002186";
         WHEN "01101110010" => data <= X"0C03319E";
         WHEN "01101110011" => data <= X"1C00619E";
         WHEN "01101110100" => data <= X"009831E2";
         WHEN "01101110101" => data <= X"00A831E2";
         WHEN "01101110110" => data <= X"0005F1DB";
         WHEN "01101110111" => data <= X"01005A9F";
         WHEN "01101111000" => data <= X"FF0020AA";
         WHEN "01101111001" => data <= X"0088BAE5";
         WHEN "01101111010" => data <= X"B7FFFF0F";
         WHEN "01101111011" => data <= X"00000015";
         WHEN "01101111100" => data <= X"B6FEFF07";
         WHEN "01101111101" => data <= X"00000015";
         WHEN "01101111110" => data <= X"E0FFFF03";
         WHEN "01101111111" => data <= X"FF004BA4";
         WHEN "01110000000" => data <= X"2D0020AA";
         WHEN "01110000001" => data <= X"008818E4";
         WHEN "01110000010" => data <= X"0B000010";
         WHEN "01110000011" => data <= X"008858E4";
         WHEN "01110000100" => data <= X"35000010";
         WHEN "01110000101" => data <= X"3D0020AA";
         WHEN "01110000110" => data <= X"2A0020AA";
         WHEN "01110000111" => data <= X"008818E4";
         WHEN "01110001000" => data <= X"69000010";
         WHEN "01110001001" => data <= X"2B0020AA";
         WHEN "01110001010" => data <= X"008818E4";
         WHEN "01110001011" => data <= X"0700000C";
         WHEN "01110001100" => data <= X"00006019";
         WHEN "01110001101" => data <= X"A5FEFF07";
         WHEN "01110001110" => data <= X"00000015";
         WHEN "01110001111" => data <= X"180020AA";
         WHEN "01110010000" => data <= X"08886BE1";
         WHEN "01110010001" => data <= X"88886BE1";
         WHEN "01110010010" => data <= X"180020AA";
         WHEN "01110010011" => data <= X"088818E3";
         WHEN "01110010100" => data <= X"888818E3";
         WHEN "01110010101" => data <= X"FFFF40AC";
         WHEN "01110010110" => data <= X"0000201A";
         WHEN "01110010111" => data <= X"FF00E0AA";
         WHEN "01110011000" => data <= X"008871E2";
         WHEN "01110011001" => data <= X"008873E2";
         WHEN "01110011010" => data <= X"0C03739E";
         WHEN "01110011011" => data <= X"1C00A19E";
         WHEN "01110011100" => data <= X"00A873E2";
         WHEN "01110011101" => data <= X"00FD3393";
         WHEN "01110011110" => data <= X"00C039E4";
         WHEN "01110011111" => data <= X"08000010";
         WHEN "01110100000" => data <= X"00000015";
         WHEN "01110100001" => data <= X"01FD7392";
         WHEN "01110100010" => data <= X"005813E4";
         WHEN "01110100011" => data <= X"0400000C";
         WHEN "01110100100" => data <= X"00000015";
         WHEN "01110100101" => data <= X"048851E0";
         WHEN "01110100110" => data <= X"000120AA";
         WHEN "01110100111" => data <= X"0100319E";
         WHEN "01110101000" => data <= X"00B8B1E5";
         WHEN "01110101001" => data <= X"F0FFFF13";
         WHEN "01110101010" => data <= X"008871E2";
         WHEN "01110101011" => data <= X"0000201A";
         WHEN "01110101100" => data <= X"008862E5";
         WHEN "01110101101" => data <= X"0502000C";
         WHEN "01110101110" => data <= X"00F0A018";
         WHEN "01110101111" => data <= X"00F0401B";
         WHEN "01110110000" => data <= X"00F0001B";
         WHEN "01110110001" => data <= X"8E1D5A9F";
         WHEN "01110110010" => data <= X"F409189F";
         WHEN "01110110011" => data <= X"0000201A";
         WHEN "01110110100" => data <= X"008832E4";
         WHEN "01110110101" => data <= X"00020010";
         WHEN "01110110110" => data <= X"00881CE4";
         WHEN "01110110111" => data <= X"7AFFFF03";
         WHEN "01110111000" => data <= X"010040AA";
         WHEN "01110111001" => data <= X"008818E4";
         WHEN "01110111010" => data <= X"D3FFFF13";
         WHEN "01110111011" => data <= X"400020AA";
         WHEN "01110111100" => data <= X"008818E4";
         WHEN "01110111101" => data <= X"D5FFFF0F";
         WHEN "01110111110" => data <= X"00006019";
         WHEN "01110111111" => data <= X"7EFEFF07";
         WHEN "01111000000" => data <= X"200060A8";
         WHEN "01111000001" => data <= X"080020AA";
         WHEN "01111000010" => data <= X"00F0A018";
         WHEN "01111000011" => data <= X"00F06018";
         WHEN "01111000100" => data <= X"08888BE2";
         WHEN "01111000101" => data <= X"005801D4";
         WHEN "01111000110" => data <= X"0A0020AA";
         WHEN "01111000111" => data <= X"831AA59C";
         WHEN "01111001000" => data <= X"00008018";
         WHEN "01111001001" => data <= X"F409639C";
         WHEN "01111001010" => data <= X"488894E2";
         WHEN "01111001011" => data <= X"D4FDFF07";
         WHEN "01111001100" => data <= X"0458CBE2";
         WHEN "01111001101" => data <= X"0000201A";
         WHEN "01111001110" => data <= X"008814E4";
         WHEN "01111001111" => data <= X"63FFFF0F";
         WHEN "01111010000" => data <= X"270040AB";
         WHEN "01111010001" => data <= X"61FFFF03";
         WHEN "01111010010" => data <= X"0000C019";
         WHEN "01111010011" => data <= X"00F0A018";
         WHEN "01111010100" => data <= X"5F1AA59C";
         WHEN "01111010101" => data <= X"00F08018";
         WHEN "01111010110" => data <= X"8C08849C";
         WHEN "01111010111" => data <= X"00F06018";
         WHEN "01111011000" => data <= X"0E000000";
         WHEN "01111011001" => data <= X"F409639C";
         WHEN "01111011010" => data <= X"00007084";
         WHEN "01111011011" => data <= X"27FFFF07";
         WHEN "01111011100" => data <= X"00000015";
         WHEN "01111011101" => data <= X"0000201A";
         WHEN "01111011110" => data <= X"00F08018";
         WHEN "01111011111" => data <= X"00F06018";
         WHEN "01111100000" => data <= X"00880BE4";
         WHEN "01111100001" => data <= X"8C08849C";
         WHEN "01111100010" => data <= X"08000010";
         WHEN "01111100011" => data <= X"F409639C";
         WHEN "01111100100" => data <= X"00F0A018";
         WHEN "01111100101" => data <= X"A11AA59C";
         WHEN "01111100110" => data <= X"B9FDFF07";
         WHEN "01111100111" => data <= X"270040AB";
         WHEN "01111101000" => data <= X"4AFFFF03";
         WHEN "01111101001" => data <= X"00000015";
         WHEN "01111101010" => data <= X"00F0A018";
         WHEN "01111101011" => data <= X"BC1AA59C";
         WHEN "01111101100" => data <= X"B3FDFF07";
         WHEN "01111101101" => data <= X"00000015";
         WHEN "01111101110" => data <= X"30000074";
         WHEN "01111101111" => data <= X"43FFFF03";
         WHEN "01111110000" => data <= X"270040AB";
         WHEN "01111110001" => data <= X"41FEFF07";
         WHEN "01111110010" => data <= X"00000015";
         WHEN "01111110011" => data <= X"FF006BA5";
         WHEN "01111110100" => data <= X"6D0020AA";
         WHEN "01111110101" => data <= X"00880BE4";
         WHEN "01111110110" => data <= X"53010010";
         WHEN "01111110111" => data <= X"00884BE4";
         WHEN "01111111000" => data <= X"50000010";
         WHEN "01111111001" => data <= X"730020AA";
         WHEN "01111111010" => data <= X"660020AA";
         WHEN "01111111011" => data <= X"00880BE4";
         WHEN "01111111100" => data <= X"F3000010";
         WHEN "01111111101" => data <= X"00884BE4";
         WHEN "01111111110" => data <= X"32000010";
         WHEN "01111111111" => data <= X"680020AA";
         WHEN "10000000000" => data <= X"630020AA";
         WHEN "10000000001" => data <= X"00880BE4";
         WHEN "10000000010" => data <= X"AA000010";
         WHEN "10000000011" => data <= X"650020AA";
         WHEN "10000000100" => data <= X"00880BE4";
         WHEN "10000000101" => data <= X"2CFFFF0F";
         WHEN "10000000110" => data <= X"00F0401B";
         WHEN "10000000111" => data <= X"00F0001B";
         WHEN "10000001000" => data <= X"8C085A9F";
         WHEN "10000001001" => data <= X"F409189F";
         WHEN "10000001010" => data <= X"00F0A018";
         WHEN "10000001011" => data <= X"871CA59C";
         WHEN "10000001100" => data <= X"04D09AE0";
         WHEN "10000001101" => data <= X"92FDFF07";
         WHEN "10000001110" => data <= X"04C078E0";
         WHEN "10000001111" => data <= X"00F04018";
         WHEN "10000010000" => data <= X"1B1CA29C";
         WHEN "10000010001" => data <= X"0004201A";
         WHEN "10000010010" => data <= X"FFFFE0AE";
         WHEN "10000010011" => data <= X"00FC201B";
         WHEN "10000010100" => data <= X"00054018";
         WHEN "10000010101" => data <= X"00007186";
         WHEN "10000010110" => data <= X"00B813E4";
         WHEN "10000010111" => data <= X"12000010";
         WHEN "10000011000" => data <= X"00C871E2";
         WHEN "10000011001" => data <= X"009801D4";
         WHEN "10000011010" => data <= X"04D09AE0";
         WHEN "10000011011" => data <= X"04C078E0";
         WHEN "10000011100" => data <= X"20B801D4";
         WHEN "10000011101" => data <= X"1CC801D4";
         WHEN "10000011110" => data <= X"188801D4";
         WHEN "10000011111" => data <= X"0C2801D4";
         WHEN "10000100000" => data <= X"7FFDFF07";
         WHEN "10000100001" => data <= X"149801D4";
         WHEN "10000100010" => data <= X"14006186";
         WHEN "10000100011" => data <= X"6FFCFF07";
         WHEN "10000100100" => data <= X"049873E0";
         WHEN "10000100101" => data <= X"2000E186";
         WHEN "10000100110" => data <= X"1C002187";
         WHEN "10000100111" => data <= X"18002186";
         WHEN "10000101000" => data <= X"0C00A184";
         WHEN "10000101001" => data <= X"0400319E";
         WHEN "10000101010" => data <= X"001031E4";
         WHEN "10000101011" => data <= X"EAFFFF13";
         WHEN "10000101100" => data <= X"00000015";
         WHEN "10000101101" => data <= X"00F0A018";
         WHEN "10000101110" => data <= X"D6000000";
         WHEN "10000101111" => data <= X"A51CA59C";
         WHEN "10000110000" => data <= X"00880BE4";
         WHEN "10000110001" => data <= X"47000010";
         WHEN "10000110010" => data <= X"690020AA";
         WHEN "10000110011" => data <= X"00880BE4";
         WHEN "10000110100" => data <= X"FEFEFF0F";
         WHEN "10000110101" => data <= X"270040AB";
         WHEN "10000110110" => data <= X"00007084";
         WHEN "10000110111" => data <= X"CBFEFF07";
         WHEN "10000111000" => data <= X"00000015";
         WHEN "10000111001" => data <= X"0000201A";
         WHEN "10000111010" => data <= X"00880BE4";
         WHEN "10000111011" => data <= X"00F08018";
         WHEN "10000111100" => data <= X"00F06018";
         WHEN "10000111101" => data <= X"04003086";
         WHEN "10000111110" => data <= X"8C08849C";
         WHEN "10000111111" => data <= X"50000010";
         WHEN "10001000000" => data <= X"F409639C";
         WHEN "10001000001" => data <= X"00F0A018";
         WHEN "10001000010" => data <= X"048801D4";
         WHEN "10001000011" => data <= X"000001D4";
         WHEN "10001000100" => data <= X"5BFDFF07";
         WHEN "10001000101" => data <= X"021BA59C";
         WHEN "10001000110" => data <= X"ECFEFF03";
         WHEN "10001000111" => data <= X"270040AB";
         WHEN "10001001000" => data <= X"00880BE4";
         WHEN "10001001001" => data <= X"39000010";
         WHEN "10001001010" => data <= X"00884BE4";
         WHEN "10001001011" => data <= X"1F000010";
         WHEN "10001001100" => data <= X"740020AA";
         WHEN "10001001101" => data <= X"700020AA";
         WHEN "10001001110" => data <= X"00880BE4";
         WHEN "10001001111" => data <= X"37000010";
         WHEN "10001010000" => data <= X"720020AA";
         WHEN "10001010001" => data <= X"00880BE4";
         WHEN "10001010010" => data <= X"DFFEFF0F";
         WHEN "10001010011" => data <= X"0004001B";
         WHEN "10001010100" => data <= X"00007884";
         WHEN "10001010101" => data <= X"ADFEFF07";
         WHEN "10001010110" => data <= X"00000015";
         WHEN "10001010111" => data <= X"0000201A";
         WHEN "10001011000" => data <= X"00882BE4";
         WHEN "10001011001" => data <= X"EE000010";
         WHEN "10001011010" => data <= X"00F0A018";
         WHEN "10001011011" => data <= X"040038AA";
         WHEN "10001011100" => data <= X"00007186";
         WHEN "10001011101" => data <= X"020020AA";
         WHEN "10001011110" => data <= X"088873E2";
         WHEN "10001011111" => data <= X"0000201A";
         WHEN "10001100000" => data <= X"008833E4";
         WHEN "10001100001" => data <= X"E1000010";
         WHEN "10001100010" => data <= X"0088B8E2";
         WHEN "10001100011" => data <= X"00F0A018";
         WHEN "10001100100" => data <= X"00F08018";
         WHEN "10001100101" => data <= X"00F06018";
         WHEN "10001100110" => data <= X"F119A59C";
         WHEN "10001100111" => data <= X"8C08849C";
         WHEN "10001101000" => data <= X"84FFFF03";
         WHEN "10001101001" => data <= X"F409639C";
         WHEN "10001101010" => data <= X"00880BE4";
         WHEN "10001101011" => data <= X"2D000010";
         WHEN "10001101100" => data <= X"760020AA";
         WHEN "10001101101" => data <= X"00880BE4";
         WHEN "10001101110" => data <= X"C3FEFF0F";
         WHEN "10001101111" => data <= X"00F0A018";
         WHEN "10001110000" => data <= X"00F08018";
         WHEN "10001110001" => data <= X"00F06018";
         WHEN "10001110010" => data <= X"ED1AA59C";
         WHEN "10001110011" => data <= X"8C08849C";
         WHEN "10001110100" => data <= X"2BFDFF07";
         WHEN "10001110101" => data <= X"F409639C";
         WHEN "10001110110" => data <= X"BBFEFF03";
         WHEN "10001110111" => data <= X"0000C01B";
         WHEN "10001111000" => data <= X"00F0A018";
         WHEN "10001111001" => data <= X"00F06018";
         WHEN "10001111010" => data <= X"BD1CA59C";
         WHEN "10001111011" => data <= X"00008018";
         WHEN "10001111100" => data <= X"23FDFF07";
         WHEN "10001111101" => data <= X"8C08639C";
         WHEN "10001111110" => data <= X"10FEFF07";
         WHEN "10001111111" => data <= X"270040AB";
         WHEN "10010000000" => data <= X"B2FEFF03";
         WHEN "10010000001" => data <= X"00000015";
         WHEN "10010000010" => data <= X"45FCFF07";
         WHEN "10010000011" => data <= X"270040AB";
         WHEN "10010000100" => data <= X"AEFEFF03";
         WHEN "10010000101" => data <= X"00000015";
         WHEN "10010000110" => data <= X"00F0A018";
         WHEN "10010000111" => data <= X"00F08018";
         WHEN "10010001000" => data <= X"00F06018";
         WHEN "10010001001" => data <= X"D91AA59C";
         WHEN "10010001010" => data <= X"8C08849C";
         WHEN "10010001011" => data <= X"14FDFF07";
         WHEN "10010001100" => data <= X"F409639C";
         WHEN "10010001101" => data <= X"A4FEFF03";
         WHEN "10010001110" => data <= X"0100C0AB";
         WHEN "10010001111" => data <= X"020060AA";
         WHEN "10010010000" => data <= X"089831E2";
         WHEN "10010010001" => data <= X"FFFF319E";
         WHEN "10010010010" => data <= X"00F0A018";
         WHEN "10010010011" => data <= X"008801D4";
         WHEN "10010010100" => data <= X"0BFDFF07";
         WHEN "10010010101" => data <= X"161BA59C";
         WHEN "10010010110" => data <= X"9CFEFF03";
         WHEN "10010010111" => data <= X"270040AB";
         WHEN "10010011000" => data <= X"0000201A";
         WHEN "10010011001" => data <= X"00F08018";
         WHEN "10010011010" => data <= X"00F06018";
         WHEN "10010011011" => data <= X"008830E4";
         WHEN "10010011100" => data <= X"8C08849C";
         WHEN "10010011101" => data <= X"09000010";
         WHEN "10010011110" => data <= X"F409639C";
         WHEN "10010011111" => data <= X"00F0A018";
         WHEN "10010100000" => data <= X"FFFCFF07";
         WHEN "10010100001" => data <= X"3F1BA59C";
         WHEN "10010100010" => data <= X"0000C019";
         WHEN "10010100011" => data <= X"0004001A";
         WHEN "10010100100" => data <= X"8EFEFF03";
         WHEN "10010100101" => data <= X"270040AB";
         WHEN "10010100110" => data <= X"00F0A018";
         WHEN "10010100111" => data <= X"F8FCFF07";
         WHEN "10010101000" => data <= X"521BA59C";
         WHEN "10010101001" => data <= X"0000C019";
         WHEN "10010101010" => data <= X"87FEFF03";
         WHEN "10010101011" => data <= X"0000001A";
         WHEN "10010101100" => data <= X"0000201A";
         WHEN "10010101101" => data <= X"008810E4";
         WHEN "10010101110" => data <= X"0B000010";
         WHEN "10010101111" => data <= X"00F0A018";
         WHEN "10010110000" => data <= X"00F08018";
         WHEN "10010110001" => data <= X"00F06018";
         WHEN "10010110010" => data <= X"651BA59C";
         WHEN "10010110011" => data <= X"8C08849C";
         WHEN "10010110100" => data <= X"F409639C";
         WHEN "10010110101" => data <= X"EAFCFF07";
         WHEN "10010110110" => data <= X"0004001A";
         WHEN "10010110111" => data <= X"7BFEFF03";
         WHEN "10010111000" => data <= X"270040AB";
         WHEN "10010111001" => data <= X"00007084";
         WHEN "10010111010" => data <= X"48FEFF07";
         WHEN "10010111011" => data <= X"00000015";
         WHEN "10010111100" => data <= X"0000201A";
         WHEN "10010111101" => data <= X"00880BE4";
         WHEN "10010111110" => data <= X"05000010";
         WHEN "10010111111" => data <= X"3F00201A";
         WHEN "10011000000" => data <= X"00F0A018";
         WHEN "10011000001" => data <= X"14FFFF03";
         WHEN "10011000010" => data <= X"871BA59C";
         WHEN "10011000011" => data <= X"FFFF31AA";
         WHEN "10011000100" => data <= X"04007086";
         WHEN "10011000101" => data <= X"0088B3E4";
         WHEN "10011000110" => data <= X"21000010";
         WHEN "10011000111" => data <= X"00F0A018";
         WHEN "10011001000" => data <= X"0DFFFF03";
         WHEN "10011001001" => data <= X"A41BA59C";
         WHEN "10011001010" => data <= X"0088B8E2";
         WHEN "10011001011" => data <= X"00007587";
         WHEN "10011001100" => data <= X"00003887";
         WHEN "10011001101" => data <= X"00C81BE4";
         WHEN "10011001110" => data <= X"10000010";
         WHEN "10011001111" => data <= X"048838E2";
         WHEN "10011010000" => data <= X"00F06018";
         WHEN "10011010001" => data <= X"0000B586";
         WHEN "10011010010" => data <= X"04D0BAE0";
         WHEN "10011010011" => data <= X"00003887";
         WHEN "10011010100" => data <= X"041082E0";
         WHEN "10011010101" => data <= X"08C801D4";
         WHEN "10011010110" => data <= X"04A801D4";
         WHEN "10011010111" => data <= X"008801D4";
         WHEN "10011011000" => data <= X"F409639C";
         WHEN "10011011001" => data <= X"14B801D4";
         WHEN "10011011010" => data <= X"C5FCFF07";
         WHEN "10011011011" => data <= X"0C9801D4";
         WHEN "10011011100" => data <= X"1400E186";
         WHEN "10011011101" => data <= X"0C006186";
         WHEN "10011011110" => data <= X"0100739E";
         WHEN "10011011111" => data <= X"0400189F";
         WHEN "10011100000" => data <= X"00003786";
         WHEN "10011100001" => data <= X"009851E4";
         WHEN "10011100010" => data <= X"E8FFFF13";
         WHEN "10011100011" => data <= X"0004201A";
         WHEN "10011100100" => data <= X"00F0A018";
         WHEN "10011100101" => data <= X"F0FEFF03";
         WHEN "10011100110" => data <= X"EA1BA59C";
         WHEN "10011100111" => data <= X"00F0401B";
         WHEN "10011101000" => data <= X"00F04018";
         WHEN "10011101001" => data <= X"0000001B";
         WHEN "10011101010" => data <= X"0000601A";
         WHEN "10011101011" => data <= X"0400E0AA";
         WHEN "10011101100" => data <= X"C41B5A9F";
         WHEN "10011101101" => data <= X"F3FFFF03";
         WHEN "10011101110" => data <= X"8C08429C";
         WHEN "10011101111" => data <= X"0000201A";
         WHEN "10011110000" => data <= X"00F0401B";
         WHEN "10011110001" => data <= X"00F0001B";
         WHEN "10011110010" => data <= X"008810E4";
         WHEN "10011110011" => data <= X"8C085A9F";
         WHEN "10011110100" => data <= X"07000010";
         WHEN "10011110101" => data <= X"F409189F";
         WHEN "10011110110" => data <= X"00F0A018";
         WHEN "10011110111" => data <= X"651BA59C";
         WHEN "10011111000" => data <= X"04D09AE0";
         WHEN "10011111001" => data <= X"BCFFFF03";
         WHEN "10011111010" => data <= X"04C078E0";
         WHEN "10011111011" => data <= X"00007084";
         WHEN "10011111100" => data <= X"06FEFF07";
         WHEN "10011111101" => data <= X"00000015";
         WHEN "10011111110" => data <= X"0000201A";
         WHEN "10011111111" => data <= X"00880BE4";
         WHEN "10100000000" => data <= X"07000010";
         WHEN "10100000001" => data <= X"3F00201A";
         WHEN "10100000010" => data <= X"00F0A018";
         WHEN "10100000011" => data <= X"871BA59C";
         WHEN "10100000100" => data <= X"04D09AE0";
         WHEN "10100000101" => data <= X"E1FEFF03";
         WHEN "10100000110" => data <= X"04C078E0";
         WHEN "10100000111" => data <= X"FFFF31AA";
         WHEN "10100001000" => data <= X"04007086";
         WHEN "10100001001" => data <= X"0088B3E4";
         WHEN "10100001010" => data <= X"04000010";
         WHEN "10100001011" => data <= X"00F0A018";
         WHEN "10100001100" => data <= X"F8FFFF03";
         WHEN "10100001101" => data <= X"A41BA59C";
         WHEN "10100001110" => data <= X"00F0A018";
         WHEN "10100001111" => data <= X"F81BA59C";
         WHEN "10100010000" => data <= X"04D09AE0";
         WHEN "10100010001" => data <= X"8EFCFF07";
         WHEN "10100010010" => data <= X"04C078E0";
         WHEN "10100010011" => data <= X"00F0A018";
         WHEN "10100010100" => data <= X"0004201A";
         WHEN "10100010101" => data <= X"0000601A";
         WHEN "10100010110" => data <= X"040040A8";
         WHEN "10100010111" => data <= X"FFFFE0AE";
         WHEN "10100011000" => data <= X"00FC201B";
         WHEN "10100011001" => data <= X"1B1CA59C";
         WHEN "10100011010" => data <= X"0000A286";
         WHEN "10100011011" => data <= X"009855E4";
         WHEN "10100011100" => data <= X"0D000010";
         WHEN "10100011101" => data <= X"04D09AE0";
         WHEN "10100011110" => data <= X"00F0A018";
         WHEN "10100011111" => data <= X"421CA59C";
         WHEN "10100100000" => data <= X"7FFCFF07";
         WHEN "10100100001" => data <= X"04C078E0";
         WHEN "10100100010" => data <= X"00006018";
         WHEN "10100100011" => data <= X"00008284";
         WHEN "10100100100" => data <= X"75FBFF07";
         WHEN "10100100101" => data <= X"00000015";
         WHEN "10100100110" => data <= X"00F0A018";
         WHEN "10100100111" => data <= X"DDFFFF03";
         WHEN "10100101000" => data <= X"5B1CA59C";
         WHEN "10100101001" => data <= X"0000B186";
         WHEN "10100101010" => data <= X"00B815E4";
         WHEN "10100101011" => data <= X"14000010";
         WHEN "10100101100" => data <= X"00C8B1E2";
         WHEN "10100101101" => data <= X"00A801D4";
         WHEN "10100101110" => data <= X"04D09AE0";
         WHEN "10100101111" => data <= X"04C078E0";
         WHEN "10100110000" => data <= X"24B801D4";
         WHEN "10100110001" => data <= X"209801D4";
         WHEN "10100110010" => data <= X"1CC801D4";
         WHEN "10100110011" => data <= X"188801D4";
         WHEN "10100110100" => data <= X"0C2801D4";
         WHEN "10100110101" => data <= X"6AFCFF07";
         WHEN "10100110110" => data <= X"14A801D4";
         WHEN "10100110111" => data <= X"1400A186";
         WHEN "10100111000" => data <= X"5AFBFF07";
         WHEN "10100111001" => data <= X"04A875E0";
         WHEN "10100111010" => data <= X"2400E186";
         WHEN "10100111011" => data <= X"20006186";
         WHEN "10100111100" => data <= X"1C002187";
         WHEN "10100111101" => data <= X"18002186";
         WHEN "10100111110" => data <= X"0C00A184";
         WHEN "10100111111" => data <= X"0100739E";
         WHEN "10101000000" => data <= X"DAFFFF03";
         WHEN "10101000001" => data <= X"0400319E";
         WHEN "10101000010" => data <= X"0000B586";
         WHEN "10101000011" => data <= X"0400319E";
         WHEN "10101000100" => data <= X"FCAFF1D7";
         WHEN "10101000101" => data <= X"1CFFFF03";
         WHEN "10101000110" => data <= X"008833E4";
         WHEN "10101000111" => data <= X"8EFEFF03";
         WHEN "10101001000" => data <= X"711CA59C";
         WHEN "10101001001" => data <= X"00F0401B";
         WHEN "10101001010" => data <= X"00F0001B";
         WHEN "10101001011" => data <= X"8C085A9F";
         WHEN "10101001100" => data <= X"F409189F";
         WHEN "10101001101" => data <= X"00F0A018";
         WHEN "10101001110" => data <= X"C01CA59C";
         WHEN "10101001111" => data <= X"04D09AE0";
         WHEN "10101010000" => data <= X"4FFCFF07";
         WHEN "10101010001" => data <= X"04C078E0";
         WHEN "10101010010" => data <= X"00F0C019";
         WHEN "10101010011" => data <= X"E21C2E9E";
         WHEN "10101010100" => data <= X"00004018";
         WHEN "10101010101" => data <= X"0C8801D4";
         WHEN "10101010110" => data <= X"04D09AE0";
         WHEN "10101010111" => data <= X"04C078E0";
         WHEN "10101011000" => data <= X"47FCFF07";
         WHEN "10101011001" => data <= X"0C00A184";
         WHEN "10101011010" => data <= X"0000201A";
         WHEN "10101011011" => data <= X"0002601A";
         WHEN "10101011100" => data <= X"0200A0AA";
         WHEN "10101011101" => data <= X"00A802E4";
         WHEN "10101011110" => data <= X"03000010";
         WHEN "10101011111" => data <= X"00000015";
         WHEN "10101100000" => data <= X"0100F172";
         WHEN "10101100001" => data <= X"008811D4";
         WHEN "10101100010" => data <= X"0400319E";
         WHEN "10101100011" => data <= X"009831E4";
         WHEN "10101100100" => data <= X"F9FFFF13";
         WHEN "10101100101" => data <= X"0200A0AA";
         WHEN "10101100110" => data <= X"00F0A018";
         WHEN "10101100111" => data <= X"EE1CA59C";
         WHEN "10101101000" => data <= X"04D09AE0";
         WHEN "10101101001" => data <= X"36FCFF07";
         WHEN "10101101010" => data <= X"04C078E0";
         WHEN "10101101011" => data <= X"0000201A";
         WHEN "10101101100" => data <= X"0000C019";
         WHEN "10101101101" => data <= X"1D0020AB";
         WHEN "10101101110" => data <= X"0002E01A";
         WHEN "10101101111" => data <= X"020060AA";
         WHEN "10101110000" => data <= X"009802E4";
         WHEN "10101110001" => data <= X"03000010";
         WHEN "10101110010" => data <= X"00000015";
         WHEN "10101110011" => data <= X"01007173";
         WHEN "10101110100" => data <= X"00007187";
         WHEN "10101110101" => data <= X"00881BE4";
         WHEN "10101110110" => data <= X"13000010";
         WHEN "10101110111" => data <= X"00C84EE4";
         WHEN "10101111000" => data <= X"10000010";
         WHEN "10101111001" => data <= X"00000015";
         WHEN "10101111010" => data <= X"00007187";
         WHEN "10101111011" => data <= X"04D09AE0";
         WHEN "10101111100" => data <= X"088801D4";
         WHEN "10101111101" => data <= X"008801D4";
         WHEN "10101111110" => data <= X"04D801D4";
         WHEN "10101111111" => data <= X"04C078E0";
         WHEN "10110000000" => data <= X"1CC801D4";
         WHEN "10110000001" => data <= X"18B801D4";
         WHEN "10110000010" => data <= X"148801D4";
         WHEN "10110000011" => data <= X"1CFCFF07";
         WHEN "10110000100" => data <= X"1000A184";
         WHEN "10110000101" => data <= X"1C002187";
         WHEN "10110000110" => data <= X"1800E186";
         WHEN "10110000111" => data <= X"14002186";
         WHEN "10110001000" => data <= X"0100CE9D";
         WHEN "10110001001" => data <= X"0400319E";
         WHEN "10110001010" => data <= X"00B831E4";
         WHEN "10110001011" => data <= X"E5FFFF13";
         WHEN "10110001100" => data <= X"020060AA";
         WHEN "10110001101" => data <= X"0000201A";
         WHEN "10110001110" => data <= X"00880EE4";
         WHEN "10110001111" => data <= X"10000010";
         WHEN "10110010000" => data <= X"030020AA";
         WHEN "10110010001" => data <= X"00F0A018";
         WHEN "10110010010" => data <= X"007001D4";
         WHEN "10110010011" => data <= X"181DA59C";
         WHEN "10110010100" => data <= X"04D09AE0";
         WHEN "10110010101" => data <= X"0AFCFF07";
         WHEN "10110010110" => data <= X"04C078E0";
         WHEN "10110010111" => data <= X"00F0A018";
         WHEN "10110011000" => data <= X"007001D4";
         WHEN "10110011001" => data <= X"311DA59C";
         WHEN "10110011010" => data <= X"04D09AE0";
         WHEN "10110011011" => data <= X"04FCFF07";
         WHEN "10110011100" => data <= X"04C078E0";
         WHEN "10110011101" => data <= X"94FDFF03";
         WHEN "10110011110" => data <= X"0000C019";
         WHEN "10110011111" => data <= X"0100429C";
         WHEN "10110100000" => data <= X"008822E4";
         WHEN "10110100001" => data <= X"B6FFFF13";
         WHEN "10110100010" => data <= X"04D09AE0";
         WHEN "10110100011" => data <= X"F5FFFF03";
         WHEN "10110100100" => data <= X"00F0A018";
         WHEN "10110100101" => data <= X"8DFCFF07";
         WHEN "10110100110" => data <= X"270040AB";
         WHEN "10110100111" => data <= X"8BFCFF07";
         WHEN "10110101000" => data <= X"FF000BA7";
         WHEN "10110101001" => data <= X"D0FF189F";
         WHEN "10110101010" => data <= X"020020AA";
         WHEN "10110101011" => data <= X"088838E2";
         WHEN "10110101100" => data <= X"FF004BA6";
         WHEN "10110101101" => data <= X"00C031E2";
         WHEN "10110101110" => data <= X"008831E2";
         WHEN "10110101111" => data <= X"D0FF529E";
         WHEN "10110110000" => data <= X"82FDFF03";
         WHEN "10110110001" => data <= X"008852E2";
         WHEN "10110110010" => data <= X"4C1DA59C";
         WHEN "10110110011" => data <= X"24FEFF03";
         WHEN "10110110100" => data <= X"00008018";
         WHEN "10110110101" => data <= X"18000010";
         WHEN "10110110110" => data <= X"080020AA";
         WHEN "10110110111" => data <= X"0888D6E2";
         WHEN "10110111000" => data <= X"01009C9F";
         WHEN "10110111001" => data <= X"040020AA";
         WHEN "10110111010" => data <= X"00883CE4";
         WHEN "10110111011" => data <= X"30000010";
         WHEN "10110111100" => data <= X"00B0C2E2";
         WHEN "10110111101" => data <= X"0000201A";
         WHEN "10110111110" => data <= X"008810E4";
         WHEN "10110111111" => data <= X"10000010";
         WHEN "10111000000" => data <= X"0000601A";
         WHEN "10111000001" => data <= X"008834E4";
         WHEN "10111000010" => data <= X"6FFDFF13";
         WHEN "10111000011" => data <= X"010040AA";
         WHEN "10111000100" => data <= X"00F0A018";
         WHEN "10111000101" => data <= X"00F08018";
         WHEN "10111000110" => data <= X"00F06018";
         WHEN "10111000111" => data <= X"5A1DA59C";
         WHEN "10111001000" => data <= X"8C08849C";
         WHEN "10111001001" => data <= X"D6FBFF07";
         WHEN "10111001010" => data <= X"F409639C";
         WHEN "10111001011" => data <= X"66FDFF03";
         WHEN "10111001100" => data <= X"049092E2";
         WHEN "10111001101" => data <= X"EBFFFF03";
         WHEN "10111001110" => data <= X"0000C01A";
         WHEN "10111001111" => data <= X"020020AA";
         WHEN "10111010000" => data <= X"088894E3";
         WHEN "10111010001" => data <= X"FF3F34A6";
         WHEN "10111010010" => data <= X"009831E4";
         WHEN "10111010011" => data <= X"07000010";
         WHEN "10111010100" => data <= X"00F0A018";
         WHEN "10111010101" => data <= X"00E001D4";
         WHEN "10111010110" => data <= X"7B1DA59C";
         WHEN "10111010111" => data <= X"00008018";
         WHEN "10111011000" => data <= X"C7FBFF07";
         WHEN "10111011001" => data <= X"04C078E0";
         WHEN "10111011010" => data <= X"0000201A";
         WHEN "10111011011" => data <= X"00881EE4";
         WHEN "10111011100" => data <= X"11000010";
         WHEN "10111011101" => data <= X"00E030E2";
         WHEN "10111011110" => data <= X"01007672";
         WHEN "10111011111" => data <= X"009811D4";
         WHEN "10111100000" => data <= X"0100949E";
         WHEN "10111100001" => data <= X"00A06EE4";
         WHEN "10111100010" => data <= X"09000010";
         WHEN "10111100011" => data <= X"0000801B";
         WHEN "10111100100" => data <= X"0000201A";
         WHEN "10111100101" => data <= X"00881EE4";
         WHEN "10111100110" => data <= X"05000010";
         WHEN "10111100111" => data <= X"00000015";
         WHEN "10111101000" => data <= X"04A010D4";
         WHEN "10111101001" => data <= X"04A0D4E1";
         WHEN "10111101010" => data <= X"0000801B";
         WHEN "10111101011" => data <= X"C8FDFF03";
         WHEN "10111101100" => data <= X"FFFF529E";
         WHEN "10111101101" => data <= X"00003186";
         WHEN "10111101110" => data <= X"01003172";
         WHEN "10111101111" => data <= X"008816E4";
         WHEN "10111110000" => data <= X"F0FFFF13";
         WHEN "10111110001" => data <= X"04D0BAE0";
         WHEN "10111110010" => data <= X"08B001D4";
         WHEN "10111110011" => data <= X"048801D4";
         WHEN "10111110100" => data <= X"00E001D4";
         WHEN "10111110101" => data <= X"00008018";
         WHEN "10111110110" => data <= X"A9FBFF07";
         WHEN "10111110111" => data <= X"04C078E0";
         WHEN "10111111000" => data <= X"E9FFFF03";
         WHEN "10111111001" => data <= X"0100949E";
         WHEN "10111111010" => data <= X"000004E4";
         WHEN "10111111011" => data <= X"000060A9";
         WHEN "10111111100" => data <= X"15000010";
         WHEN "10111111101" => data <= X"000083A9";
         WHEN "10111111110" => data <= X"0100C0A8";
         WHEN "10111111111" => data <= X"000084E5";
         WHEN "11000000000" => data <= X"05000010";
         WHEN "11000000001" => data <= X"006084E4";
         WHEN "11000000010" => data <= X"002084E0";
         WHEN "11000000011" => data <= X"FCFFFF13";
         WHEN "11000000100" => data <= X"0030C6E0";
         WHEN "11000000101" => data <= X"0030EBE0";
         WHEN "11000000110" => data <= X"4100C6B8";
         WHEN "11000000111" => data <= X"02200CE1";
         WHEN "11000001000" => data <= X"0060A4E4";
         WHEN "11000001001" => data <= X"410084B8";
         WHEN "11000001010" => data <= X"0400000C";
         WHEN "11000001011" => data <= X"00000015";
         WHEN "11000001100" => data <= X"000067A9";
         WHEN "11000001101" => data <= X"000088A9";
         WHEN "11000001110" => data <= X"000026E4";
         WHEN "11000001111" => data <= X"F7FFFF13";
         WHEN "11000010000" => data <= X"0030EBE0";
         WHEN "11000010001" => data <= X"00480044";
         WHEN "11000010010" => data <= X"00000015";
         WHEN "11000010011" => data <= X"0000A9A9";
         WHEN "11000010100" => data <= X"E6FFFF07";
         WHEN "11000010101" => data <= X"00000015";
         WHEN "11000010110" => data <= X"00680044";
         WHEN "11000010111" => data <= X"00006CA9";
         WHEN "11000011000" => data <= X"65202449";
         WHEN "11000011001" => data <= X"726F7272";
         WHEN "11000011010" => data <= X"44000A21";
         WHEN "11000011011" => data <= X"72652024";
         WHEN "11000011100" => data <= X"0A726F72";
         WHEN "11000011101" => data <= X"71726900";
         WHEN "11000011110" => data <= X"3F3F000A";
         WHEN "11000011111" => data <= X"73000A3F";
         WHEN "11000100000" => data <= X"65747379";
         WHEN "11000100001" => data <= X"000A216D";
         WHEN "11000100010" => data <= X"63656843";
         WHEN "11000100011" => data <= X"676E696B";
         WHEN "11000100100" => data <= X"73616C20";
         WHEN "11000100101" => data <= X"61702074";
         WHEN "11000100110" => data <= X"6F206567";
         WHEN "11000100111" => data <= X"6C662066";
         WHEN "11000101000" => data <= X"20687361";
         WHEN "11000101001" => data <= X"74706D65";
         WHEN "11000101010" => data <= X"46000A79";
         WHEN "11000101011" => data <= X"6873616C";
         WHEN "11000101100" => data <= X"72726520";
         WHEN "11000101101" => data <= X"0A21726F";
         WHEN "11000101110" => data <= X"61724500";
         WHEN "11000101111" => data <= X"676E6973";
         WHEN "11000110000" => data <= X"73616C20";
         WHEN "11000110001" => data <= X"61702074";
         WHEN "11000110010" => data <= X"6F206567";
         WHEN "11000110011" => data <= X"6C462066";
         WHEN "11000110100" => data <= X"0A687361";
         WHEN "11000110101" => data <= X"69725700";
         WHEN "11000110110" => data <= X"676E6974";
         WHEN "11000110111" => data <= X"73657420";
         WHEN "11000111000" => data <= X"65732074";
         WHEN "11000111001" => data <= X"6E657571";
         WHEN "11000111010" => data <= X"74206563";
         WHEN "11000111011" => data <= X"6C66206F";
         WHEN "11000111100" => data <= X"2E687361";
         WHEN "11000111101" => data <= X"6556000A";
         WHEN "11000111110" => data <= X"79666972";
         WHEN "11000111111" => data <= X"20676E69";
         WHEN "11001000000" => data <= X"74736574";
         WHEN "11001000001" => data <= X"71657320";
         WHEN "11001000010" => data <= X"636E6575";
         WHEN "11001000011" => data <= X"72662065";
         WHEN "11001000100" => data <= X"66206D6F";
         WHEN "11001000101" => data <= X"6873616C";
         WHEN "11001000110" => data <= X"54000A2E";
         WHEN "11001000111" => data <= X"20747365";
         WHEN "11001001000" => data <= X"6C696166";
         WHEN "11001001001" => data <= X"203A6465";
         WHEN "11001001010" => data <= X"3A206425";
         WHEN "11001001011" => data <= X"25783020";
         WHEN "11001001100" => data <= X"3D2F2058";
         WHEN "11001001101" => data <= X"25783020";
         WHEN "11001001110" => data <= X"46000A58";
         WHEN "11001001111" => data <= X"6873616C";
         WHEN "11001010000" => data <= X"73657420";
         WHEN "11001010001" => data <= X"6B6F2074";
         WHEN "11001010010" => data <= X"0A2E7961";
         WHEN "11001010011" => data <= X"5343000A";
         WHEN "11001010100" => data <= X"3637342D";
         WHEN "11001010101" => data <= X"626D4520";
         WHEN "11001010110" => data <= X"65646465";
         WHEN "11001010111" => data <= X"79532064";
         WHEN "11001011000" => data <= X"6D657473";
         WHEN "11001011001" => data <= X"73654420";
         WHEN "11001011010" => data <= X"0A6E6769";
         WHEN "11001011011" => data <= X"65704F00";
         WHEN "11001011100" => data <= X"7369726E";
         WHEN "11001011101" => data <= X"61622063";
         WHEN "11001011110" => data <= X"20646573";
         WHEN "11001011111" => data <= X"74726976";
         WHEN "11001100000" => data <= X"206C6175";
         WHEN "11001100001" => data <= X"746F7250";
         WHEN "11001100010" => data <= X"7079746F";
         WHEN "11001100011" => data <= X"000A2E65";
         WHEN "11001100100" => data <= X"6C697542";
         WHEN "11001100101" => data <= X"65762064";
         WHEN "11001100110" => data <= X"6F697372";
         WHEN "11001100111" => data <= X"4D203A6E";
         WHEN "11001101000" => data <= X"53206E6F";
         WHEN "11001101001" => data <= X"20207065";
         WHEN "11001101010" => data <= X"31312032";
         WHEN "11001101011" => data <= X"3A39303A";
         WHEN "11001101100" => data <= X"41203733";
         WHEN "11001101101" => data <= X"4543204D";
         WHEN "11001101110" => data <= X"32205453";
         WHEN "11001101111" => data <= X"0A343230";
         WHEN "11001110000" => data <= X"2049000A";
         WHEN "11001110001" => data <= X"43206D61";
         WHEN "11001110010" => data <= X"25205550";
         WHEN "11001110011" => data <= X"666F2064";
         WHEN "11001110100" => data <= X"20642520";
         WHEN "11001110101" => data <= X"6E6E7572";
         WHEN "11001110110" => data <= X"20676E69";
         WHEN "11001110111" => data <= X"00207461";
         WHEN "11001111000" => data <= X"64256425";
         WHEN "11001111001" => data <= X"2564252E";
         WHEN "11001111010" => data <= X"484D2064";
         WHEN "11001111011" => data <= X"0A0A2E7A";
         WHEN "11001111100" => data <= X"65784500";
         WHEN "11001111101" => data <= X"69747563";
         WHEN "11001111110" => data <= X"6620676E";
         WHEN "11001111111" => data <= X"6873616C";
         WHEN "11010000000" => data <= X"6F727020";
         WHEN "11010000001" => data <= X"6D617267";
         WHEN "11010000010" => data <= X"0A2E2E2E";
         WHEN "11010000011" => data <= X"6F725000";
         WHEN "11010000100" => data <= X"6D617267";
         WHEN "11010000101" => data <= X"65727020";
         WHEN "11010000110" => data <= X"746E6573";
         WHEN "11010000111" => data <= X"74756220";
         WHEN "11010001000" => data <= X"746F6E20";
         WHEN "11010001001" => data <= X"726F6620";
         WHEN "11010001010" => data <= X"69687420";
         WHEN "11010001011" => data <= X"61542073";
         WHEN "11010001100" => data <= X"74656772";
         WHEN "11010001101" => data <= X"69440A2E";
         WHEN "11010001110" => data <= X"6F792064";
         WHEN "11010001111" => data <= X"70752075";
         WHEN "11010010000" => data <= X"64616F6C";
         WHEN "11010010001" => data <= X"726F6620";
         WHEN "11010010010" => data <= X"65687420";
         WHEN "11010010011" => data <= X"31524F20";
         WHEN "11010010100" => data <= X"20303234";
         WHEN "11010010101" => data <= X"74616C70";
         WHEN "11010010110" => data <= X"6D726F66";
         WHEN "11010010111" => data <= X"44000A3F";
         WHEN "11010011000" => data <= X"6C6E776F";
         WHEN "11010011001" => data <= X"3A64616F";
         WHEN "11010011010" => data <= X"6E6F6420";
         WHEN "11010011011" => data <= X"52000A65";
         WHEN "11010011100" => data <= X"69646165";
         WHEN "11010011101" => data <= X"6320676E";
         WHEN "11010011110" => data <= X"2065646F";
         WHEN "11010011111" => data <= X"6C626174";
         WHEN "11010100000" => data <= X"44000A65";
         WHEN "11010100001" => data <= X"6C6E776F";
         WHEN "11010100010" => data <= X"3A64616F";
         WHEN "11010100011" => data <= X"74657320";
         WHEN "11010100100" => data <= X"64646120";
         WHEN "11010100101" => data <= X"73736572";
         WHEN "11010100110" => data <= X"30203D20";
         WHEN "11010100111" => data <= X"0A582578";
         WHEN "11010101000" => data <= X"72724500";
         WHEN "11010101001" => data <= X"202C726F";
         WHEN "11010101010" => data <= X"70206F6E";
         WHEN "11010101011" => data <= X"72676F72";
         WHEN "11010101100" => data <= X"6C206D61";
         WHEN "11010101101" => data <= X"6564616F";
         WHEN "11010101110" => data <= X"000A2164";
         WHEN "11010101111" => data <= X"63657845";
         WHEN "11010110000" => data <= X"6E697475";
         WHEN "11010110001" => data <= X"6F6C2067";
         WHEN "11010110010" => data <= X"64656461";
         WHEN "11010110011" => data <= X"6F727020";
         WHEN "11010110100" => data <= X"6D617267";
         WHEN "11010110101" => data <= X"0A2E2E2E";
         WHEN "11010110110" => data <= X"74655300";
         WHEN "11010110111" => data <= X"676E6974";
         WHEN "11010111000" => data <= X"6F727020";
         WHEN "11010111001" => data <= X"6D202E67";
         WHEN "11010111010" => data <= X"0A65646F";
         WHEN "11010111011" => data <= X"74655300";
         WHEN "11010111100" => data <= X"676E6974";
         WHEN "11010111101" => data <= X"72657620";
         WHEN "11010111110" => data <= X"202E6669";
         WHEN "11010111111" => data <= X"65646F6D";
         WHEN "11011000000" => data <= X"6F4E000A";
         WHEN "11011000001" => data <= X"6F727020";
         WHEN "11011000010" => data <= X"6D617267";
         WHEN "11011000011" => data <= X"65727020";
         WHEN "11011000100" => data <= X"746E6573";
         WHEN "11011000101" => data <= X"7250000A";
         WHEN "11011000110" => data <= X"6172676F";
         WHEN "11011000111" => data <= X"6E69206D";
         WHEN "11011001000" => data <= X"6D656D20";
         WHEN "11011001001" => data <= X"6F726620";
         WHEN "11011001010" => data <= X"6162206D";
         WHEN "11011001011" => data <= X"302B6573";
         WHEN "11011001100" => data <= X"206F7420";
         WHEN "11011001101" => data <= X"65736162";
         WHEN "11011001110" => data <= X"2578302B";
         WHEN "11011001111" => data <= X"53000A58";
         WHEN "11011010000" => data <= X"63746977";
         WHEN "11011010001" => data <= X"20646568";
         WHEN "11011010010" => data <= X"46206F74";
         WHEN "11011010011" => data <= X"6873616C";
         WHEN "11011010100" => data <= X"7753000A";
         WHEN "11011010101" => data <= X"68637469";
         WHEN "11011010110" => data <= X"74206465";
         WHEN "11011010111" => data <= X"4453206F";
         WHEN "11011011000" => data <= X"0A6D6152";
         WHEN "11011011001" => data <= X"656C5000";
         WHEN "11011011010" => data <= X"20657361";
         WHEN "11011011011" => data <= X"6E616863";
         WHEN "11011011100" => data <= X"74206567";
         WHEN "11011011101" => data <= X"6874206F";
         WHEN "11011011110" => data <= X"44532065";
         WHEN "11011011111" => data <= X"204D4152";
         WHEN "11011100000" => data <= X"2A207962";
         WHEN "11011100001" => data <= X"4E000A74";
         WHEN "11011100010" => data <= X"7270206F";
         WHEN "11011100011" => data <= X"6172676F";
         WHEN "11011100100" => data <= X"6F6C206D";
         WHEN "11011100101" => data <= X"64656461";
         WHEN "11011100110" => data <= X"206E6920";
         WHEN "11011100111" => data <= X"61524453";
         WHEN "11011101000" => data <= X"000A216D";
         WHEN "11011101001" => data <= X"676F7250";
         WHEN "11011101010" => data <= X"206D6172";
         WHEN "11011101011" => data <= X"73656F64";
         WHEN "11011101100" => data <= X"746F6E20";
         WHEN "11011101101" => data <= X"74696620";
         WHEN "11011101110" => data <= X"206E6920";
         WHEN "11011101111" => data <= X"73616C46";
         WHEN "11011110000" => data <= X"000A2168";
         WHEN "11011110001" => data <= X"706D6F43";
         WHEN "11011110010" => data <= X"20657261";
         WHEN "11011110011" => data <= X"6F727265";
         WHEN "11011110100" => data <= X"74612072";
         WHEN "11011110101" => data <= X"25783020";
         WHEN "11011110110" => data <= X"203A2058";
         WHEN "11011110111" => data <= X"58257830";
         WHEN "11011111000" => data <= X"203D2120";
         WHEN "11011111001" => data <= X"58257830";
         WHEN "11011111010" => data <= X"6F43000A";
         WHEN "11011111011" => data <= X"7261706D";
         WHEN "11011111100" => data <= X"6F642065";
         WHEN "11011111101" => data <= X"000A656E";
         WHEN "11011111110" => data <= X"63656843";
         WHEN "11011111111" => data <= X"676E696B";
         WHEN "11100000000" => data <= X"20666920";
         WHEN "11100000001" => data <= X"20656874";
         WHEN "11100000010" => data <= X"73616C66";
         WHEN "11100000011" => data <= X"73692068";
         WHEN "11100000100" => data <= X"706D6520";
         WHEN "11100000101" => data <= X"2E2E7974";
         WHEN "11100000110" => data <= X"53000A2E";
         WHEN "11100000111" => data <= X"74726174";
         WHEN "11100001000" => data <= X"616C6620";
         WHEN "11100001001" => data <= X"65206873";
         WHEN "11100001010" => data <= X"65736172";
         WHEN "11100001011" => data <= X"63796320";
         WHEN "11100001100" => data <= X"6620656C";
         WHEN "11100001101" => data <= X"7020726F";
         WHEN "11100001110" => data <= X"20656761";
         WHEN "11100001111" => data <= X"58257830";
         WHEN "11100010000" => data <= X"7453000A";
         WHEN "11100010001" => data <= X"20747261";
         WHEN "11100010010" => data <= X"676F7270";
         WHEN "11100010011" => data <= X"6D6D6172";
         WHEN "11100010100" => data <= X"20676E69";
         WHEN "11100010101" => data <= X"73616C66";
         WHEN "11100010110" => data <= X"50000A68";
         WHEN "11100010111" => data <= X"72676F72";
         WHEN "11100011000" => data <= X"696D6D61";
         WHEN "11100011001" => data <= X"6620676E";
         WHEN "11100011010" => data <= X"73696E69";
         WHEN "11100011011" => data <= X"0A646568";
         WHEN "11100011100" => data <= X"206F4E00";
         WHEN "11100011101" => data <= X"676F7270";
         WHEN "11100011110" => data <= X"206D6172";
         WHEN "11100011111" => data <= X"66206E69";
         WHEN "11100100000" => data <= X"6873616C";
         WHEN "11100100001" => data <= X"43000A21";
         WHEN "11100100010" => data <= X"6B636568";
         WHEN "11100100011" => data <= X"20676E69";
         WHEN "11100100100" => data <= X"66206669";
         WHEN "11100100101" => data <= X"6873616C";
         WHEN "11100100110" => data <= X"20736920";
         WHEN "11100100111" => data <= X"72696427";
         WHEN "11100101000" => data <= X"0A277974";
         WHEN "11100101001" => data <= X"616C4600";
         WHEN "11100101010" => data <= X"69206873";
         WHEN "11100101011" => data <= X"6D652073";
         WHEN "11100101100" => data <= X"20797470";
         WHEN "11100101101" => data <= X"61726528";
         WHEN "11100101110" => data <= X"29646573";
         WHEN "11100101111" => data <= X"000A0A2E";
         WHEN "11100110000" => data <= X"72617453";
         WHEN "11100110001" => data <= X"676E6974";
         WHEN "11100110010" => data <= X"6D697320";
         WHEN "11100110011" => data <= X"20656C70";
         WHEN "11100110100" => data <= X"61524453";
         WHEN "11100110101" => data <= X"656D206D";
         WHEN "11100110110" => data <= X"6568636D";
         WHEN "11100110111" => data <= X"0A2E6B63";
         WHEN "11100111000" => data <= X"7257000A";
         WHEN "11100111001" => data <= X"6E697469";
         WHEN "11100111010" => data <= X"2E2E2E67";
         WHEN "11100111011" => data <= X"6556000A";
         WHEN "11100111100" => data <= X"79666972";
         WHEN "11100111101" => data <= X"2E676E69";
         WHEN "11100111110" => data <= X"000A2E2E";
         WHEN "11100111111" => data <= X"6F727245";
         WHEN "11101000000" => data <= X"30402072";
         WHEN "11101000001" => data <= X"20582578";
         WHEN "11101000010" => data <= X"7830203A";
         WHEN "11101000011" => data <= X"21205825";
         WHEN "11101000100" => data <= X"7830203D";
         WHEN "11101000101" => data <= X"000A5825";
         WHEN "11101000110" => data <= X"6F20724E";
         WHEN "11101000111" => data <= X"72652066";
         WHEN "11101001000" => data <= X"73726F72";
         WHEN "11101001001" => data <= X"756F6620";
         WHEN "11101001010" => data <= X"3A20646E";
         WHEN "11101001011" => data <= X"0A642520";
         WHEN "11101001100" => data <= X"6D654D00";
         WHEN "11101001101" => data <= X"63656863";
         WHEN "11101001110" => data <= X"6F64206B";
         WHEN "11101001111" => data <= X"202C656E";
         WHEN "11101010000" => data <= X"65206425";
         WHEN "11101010001" => data <= X"726F7272";
         WHEN "11101010010" => data <= X"000A0A73";
         WHEN "11101010011" => data <= X"6E6B6E55";
         WHEN "11101010100" => data <= X"206E776F";
         WHEN "11101010101" => data <= X"65646F63";
         WHEN "11101010110" => data <= X"61430021";
         WHEN "11101010111" => data <= X"746F6E6E";
         WHEN "11101011000" => data <= X"6F727020";
         WHEN "11101011001" => data <= X"6D617267";
         WHEN "11101011010" => data <= X"616C6620";
         WHEN "11101011011" => data <= X"202C6873";
         WHEN "11101011100" => data <= X"726F6261";
         WHEN "11101011101" => data <= X"676E6974";
         WHEN "11101011110" => data <= X"44000A21";
         WHEN "11101011111" => data <= X"6C6E776F";
         WHEN "11101100000" => data <= X"3A64616F";
         WHEN "11101100001" => data <= X"20746120";
         WHEN "11101100010" => data <= X"58257830";
         WHEN "11101100011" => data <= X"6556000A";
         WHEN "11101100100" => data <= X"69666972";
         WHEN "11101100101" => data <= X"69746163";
         WHEN "11101100110" => data <= X"65206E6F";
         WHEN "11101100111" => data <= X"726F7272";
         WHEN "11101101000" => data <= X"20746120";
         WHEN "11101101001" => data <= X"58257830";
         WHEN "11101101010" => data <= X"30203A20";
         WHEN "11101101011" => data <= X"20582578";
         WHEN "11101101100" => data <= X"30203D21";
         WHEN "11101101101" => data <= X"0A582578";
         WHEN "11101101110" => data <= X"6F6E4B00";
         WHEN "11101101111" => data <= X"52206E77";
         WHEN "11101110000" => data <= X"32333253";
         WHEN "11101110001" => data <= X"6D6F6320";
         WHEN "11101110010" => data <= X"646E616D";
         WHEN "11101110011" => data <= X"000A3A73";
         WHEN "11101110100" => data <= X"53202024";
         WHEN "11101110101" => data <= X"74726174";
         WHEN "11101110110" => data <= X"65687420";
         WHEN "11101110111" => data <= X"6F727020";
         WHEN "11101111000" => data <= X"6D617267";
         WHEN "11101111001" => data <= X"616F6C20";
         WHEN "11101111010" => data <= X"20646564";
         WHEN "11101111011" => data <= X"74206E69";
         WHEN "11101111100" => data <= X"65677261";
         WHEN "11101111101" => data <= X"2A000A74";
         WHEN "11101111110" => data <= X"65532070";
         WHEN "11101111111" => data <= X"72702074";
         WHEN "11110000000" => data <= X"6172676F";
         WHEN "11110000001" => data <= X"6E696D6D";
         WHEN "11110000010" => data <= X"6F6D2067";
         WHEN "11110000011" => data <= X"28206564";
         WHEN "11110000100" => data <= X"61666564";
         WHEN "11110000101" => data <= X"29746C75";
         WHEN "11110000110" => data <= X"762A000A";
         WHEN "11110000111" => data <= X"74655320";
         WHEN "11110001000" => data <= X"72657620";
         WHEN "11110001001" => data <= X"63696669";
         WHEN "11110001010" => data <= X"6F697461";
         WHEN "11110001011" => data <= X"6F6D206E";
         WHEN "11110001100" => data <= X"000A6564";
         WHEN "11110001101" => data <= X"5320692A";
         WHEN "11110001110" => data <= X"20776F68";
         WHEN "11110001111" => data <= X"6F666E69";
         WHEN "11110010000" => data <= X"206E6F20";
         WHEN "11110010001" => data <= X"676F7270";
         WHEN "11110010010" => data <= X"206D6172";
         WHEN "11110010011" => data <= X"74206E69";
         WHEN "11110010100" => data <= X"65677261";
         WHEN "11110010101" => data <= X"2A000A74";
         WHEN "11110010110" => data <= X"6F542074";
         WHEN "11110010111" => data <= X"656C6767";
         WHEN "11110011000" => data <= X"72617420";
         WHEN "11110011001" => data <= X"20746567";
         WHEN "11110011010" => data <= X"77746562";
         WHEN "11110011011" => data <= X"206E6565";
         WHEN "11110011100" => data <= X"61524453";
         WHEN "11110011101" => data <= X"6428206D";
         WHEN "11110011110" => data <= X"75616665";
         WHEN "11110011111" => data <= X"2029746C";
         WHEN "11110100000" => data <= X"20646E61";
         WHEN "11110100001" => data <= X"73616C46";
         WHEN "11110100010" => data <= X"2A000A68";
         WHEN "11110100011" => data <= X"6550206D";
         WHEN "11110100100" => data <= X"726F6672";
         WHEN "11110100101" => data <= X"6973206D";
         WHEN "11110100110" => data <= X"656C706D";
         WHEN "11110100111" => data <= X"52445320";
         WHEN "11110101000" => data <= X"6D206D61";
         WHEN "11110101001" => data <= X"68636D65";
         WHEN "11110101010" => data <= X"0A6B6365";
         WHEN "11110101011" => data <= X"20732A00";
         WHEN "11110101100" => data <= X"63656843";
         WHEN "11110101101" => data <= X"5053206B";
         WHEN "11110101110" => data <= X"6C662D49";
         WHEN "11110101111" => data <= X"20687361";
         WHEN "11110110000" => data <= X"70696863";
         WHEN "11110110001" => data <= X"652A000A";
         WHEN "11110110010" => data <= X"61724520";
         WHEN "11110110011" => data <= X"53206573";
         WHEN "11110110100" => data <= X"662D4950";
         WHEN "11110110101" => data <= X"6873616C";
         WHEN "11110110110" => data <= X"69686320";
         WHEN "11110110111" => data <= X"2A000A70";
         WHEN "11110111000" => data <= X"75522072";
         WHEN "11110111001" => data <= X"7270206E";
         WHEN "11110111010" => data <= X"6172676F";
         WHEN "11110111011" => data <= X"6E69206D";
         WHEN "11110111100" => data <= X"49505320";
         WHEN "11110111101" => data <= X"616C662D";
         WHEN "11110111110" => data <= X"000A6873";
         WHEN "11110111111" => data <= X"5320662A";
         WHEN "11111000000" => data <= X"65726F74";
         WHEN "11111000001" => data <= X"6F727020";
         WHEN "11111000010" => data <= X"6D617267";
         WHEN "11111000011" => data <= X"616F6C20";
         WHEN "11111000100" => data <= X"20646564";
         WHEN "11111000101" => data <= X"53206E69";
         WHEN "11111000110" => data <= X"4D415244";
         WHEN "11111000111" => data <= X"206F7420";
         WHEN "11111001000" => data <= X"2D495053";
         WHEN "11111001001" => data <= X"73616C46";
         WHEN "11111001010" => data <= X"2A000A68";
         WHEN "11111001011" => data <= X"6F432063";
         WHEN "11111001100" => data <= X"7261706D";
         WHEN "11111001101" => data <= X"72702065";
         WHEN "11111001110" => data <= X"6172676F";
         WHEN "11111001111" => data <= X"6F6C206D";
         WHEN "11111010000" => data <= X"64656461";
         WHEN "11111010001" => data <= X"206E6920";
         WHEN "11111010010" => data <= X"41524453";
         WHEN "11111010011" => data <= X"6977204D";
         WHEN "11111010100" => data <= X"53206874";
         WHEN "11111010101" => data <= X"462D4950";
         WHEN "11111010110" => data <= X"6873616C";
         WHEN "11111010111" => data <= X"682A000A";
         WHEN "11111011000" => data <= X"69685420";
         WHEN "11111011001" => data <= X"65682073";
         WHEN "11111011010" => data <= X"6373706C";
         WHEN "11111011011" => data <= X"6E656572";
         WHEN "11111011100" => data <= X"00000A0A";
         WHEN "11111011101" => data <= X"EFBEADDE";
         WHEN "11111011110" => data <= X"01000000";
         WHEN "11111011111" => data <= X"02000000";
         WHEN "11111100000" => data <= X"03000000";
         WHEN "11111100001" => data <= X"04000000";
         WHEN "11111100010" => data <= X"05000000";
         WHEN "11111100011" => data <= X"06000000";
         WHEN "11111100100" => data <= X"07000000";
         WHEN "11111100101" => data <= X"B91D00F0";
         WHEN "11111100110" => data <= X"D01D00F0";
         WHEN "11111100111" => data <= X"F71D00F0";
         WHEN "11111101000" => data <= X"1A1E00F0";
         WHEN "11111101001" => data <= X"341E00F0";
         WHEN "11111101010" => data <= X"571E00F0";
         WHEN "11111101011" => data <= X"8B1E00F0";
         WHEN "11111101100" => data <= X"AD1E00F0";
         WHEN "11111101101" => data <= X"C61E00F0";
         WHEN "11111101110" => data <= X"DF1E00F0";
         WHEN "11111101111" => data <= X"FC1E00F0";
         WHEN "11111110000" => data <= X"2B1F00F0";
         WHEN "11111110001" => data <= X"5E1F00F0";
         WHEN "11111110011" => data <= X"10000000";
         WHEN "11111110101" => data <= X"00527A01";
         WHEN "11111110110" => data <= X"01097C04";
         WHEN "11111110111" => data <= X"00010D1B";
         WHEN "11111111000" => data <= X"14000000";
         WHEN "11111111001" => data <= X"18000000";
         WHEN "11111111010" => data <= X"64F8FFFF";
         WHEN "11111111011" => data <= X"14000000";
         WHEN "11111111100" => data <= X"09094100";
         WHEN "11111111101" => data <= X"0000000D";
         WHEN OTHERS => data <= X"00000000";
      END CASE;
   END PROCESS TheRom;

END platform_independent;
